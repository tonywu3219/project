##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 10:37:00 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 570.0000 BY 470.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 284.8550 469.5300 284.9450 470.0000 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 314.9500 0.5200 315.0500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 311.9500 0.5200 312.0500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 308.9500 0.5200 309.0500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 305.9500 0.5200 306.0500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 302.9500 0.5200 303.0500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 299.9500 0.5200 300.0500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 296.9500 0.5200 297.0500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 293.9500 0.5200 294.0500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 290.9500 0.5200 291.0500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 287.9500 0.5200 288.0500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 284.9500 0.5200 285.0500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 281.9500 0.5200 282.0500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 278.9500 0.5200 279.0500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 275.9500 0.5200 276.0500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 272.9500 0.5200 273.0500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 269.9500 0.5200 270.0500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 266.9500 0.5200 267.0500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 263.9500 0.5200 264.0500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 260.9500 0.5200 261.0500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 257.9500 0.5200 258.0500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 254.9500 0.5200 255.0500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 251.9500 0.5200 252.0500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 248.9500 0.5200 249.0500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 245.9500 0.5200 246.0500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 242.9500 0.5200 243.0500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 239.9500 0.5200 240.0500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 236.9500 0.5200 237.0500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 233.9500 0.5200 234.0500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 230.9500 0.5200 231.0500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 227.9500 0.5200 228.0500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 224.9500 0.5200 225.0500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 221.9500 0.5200 222.0500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 218.9500 0.5200 219.0500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 215.9500 0.5200 216.0500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 212.9500 0.5200 213.0500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 209.9500 0.5200 210.0500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 206.9500 0.5200 207.0500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 203.9500 0.5200 204.0500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 200.9500 0.5200 201.0500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 197.9500 0.5200 198.0500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 194.9500 0.5200 195.0500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 191.9500 0.5200 192.0500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 188.9500 0.5200 189.0500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 185.9500 0.5200 186.0500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 182.9500 0.5200 183.0500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 179.9500 0.5200 180.0500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 176.9500 0.5200 177.0500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 173.9500 0.5200 174.0500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 170.9500 0.5200 171.0500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 167.9500 0.5200 168.0500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 164.9500 0.5200 165.0500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 161.9500 0.5200 162.0500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 158.9500 0.5200 159.0500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 155.9500 0.5200 156.0500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 152.9500 0.5200 153.0500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 149.9500 0.5200 150.0500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 146.9500 0.5200 147.0500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 143.9500 0.5200 144.0500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 140.9500 0.5200 141.0500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 137.9500 0.5200 138.0500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 134.9500 0.5200 135.0500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 131.9500 0.5200 132.0500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 128.9500 0.5200 129.0500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 125.9500 0.5200 126.0500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 491.4550 0.0000 491.5450 0.4700 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 488.8550 0.0000 488.9450 0.4700 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 486.2550 0.0000 486.3450 0.4700 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 483.6550 0.0000 483.7450 0.4700 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 481.0550 0.0000 481.1450 0.4700 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 478.4550 0.0000 478.5450 0.4700 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 475.8550 0.0000 475.9450 0.4700 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 473.2550 0.0000 473.3450 0.4700 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 470.6550 0.0000 470.7450 0.4700 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 468.0550 0.0000 468.1450 0.4700 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 465.4550 0.0000 465.5450 0.4700 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 462.8550 0.0000 462.9450 0.4700 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 460.2550 0.0000 460.3450 0.4700 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 457.6550 0.0000 457.7450 0.4700 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 455.0550 0.0000 455.1450 0.4700 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 452.4550 0.0000 452.5450 0.4700 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 449.8550 0.0000 449.9450 0.4700 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 447.2550 0.0000 447.3450 0.4700 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 444.6550 0.0000 444.7450 0.4700 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 442.0550 0.0000 442.1450 0.4700 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 439.4550 0.0000 439.5450 0.4700 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 436.8550 0.0000 436.9450 0.4700 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 434.2550 0.0000 434.3450 0.4700 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 431.6550 0.0000 431.7450 0.4700 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 429.0550 0.0000 429.1450 0.4700 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 426.4550 0.0000 426.5450 0.4700 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 423.8550 0.0000 423.9450 0.4700 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 421.2550 0.0000 421.3450 0.4700 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 418.6550 0.0000 418.7450 0.4700 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 416.0550 0.0000 416.1450 0.4700 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 413.4550 0.0000 413.5450 0.4700 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 410.8550 0.0000 410.9450 0.4700 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 408.2550 0.0000 408.3450 0.4700 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 405.6550 0.0000 405.7450 0.4700 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 403.0550 0.0000 403.1450 0.4700 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 400.4550 0.0000 400.5450 0.4700 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 397.8550 0.0000 397.9450 0.4700 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 395.2550 0.0000 395.3450 0.4700 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 392.6550 0.0000 392.7450 0.4700 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 390.0550 0.0000 390.1450 0.4700 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 387.4550 0.0000 387.5450 0.4700 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 384.8550 0.0000 384.9450 0.4700 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 382.2550 0.0000 382.3450 0.4700 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 379.6550 0.0000 379.7450 0.4700 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 377.0550 0.0000 377.1450 0.4700 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 374.4550 0.0000 374.5450 0.4700 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 371.8550 0.0000 371.9450 0.4700 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 369.2550 0.0000 369.3450 0.4700 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 366.6550 0.0000 366.7450 0.4700 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 364.0550 0.0000 364.1450 0.4700 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 361.4550 0.0000 361.5450 0.4700 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 358.8550 0.0000 358.9450 0.4700 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 356.2550 0.0000 356.3450 0.4700 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 353.6550 0.0000 353.7450 0.4700 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 351.0550 0.0000 351.1450 0.4700 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 348.4550 0.0000 348.5450 0.4700 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 345.8550 0.0000 345.9450 0.4700 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 343.2550 0.0000 343.3450 0.4700 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 340.6550 0.0000 340.7450 0.4700 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 338.0550 0.0000 338.1450 0.4700 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 335.4550 0.0000 335.5450 0.4700 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 332.8550 0.0000 332.9450 0.4700 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 330.2550 0.0000 330.3450 0.4700 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 327.6550 0.0000 327.7450 0.4700 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 325.0550 0.0000 325.1450 0.4700 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 322.4550 0.0000 322.5450 0.4700 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 319.8550 0.0000 319.9450 0.4700 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 317.2550 0.0000 317.3450 0.4700 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 314.6550 0.0000 314.7450 0.4700 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 312.0550 0.0000 312.1450 0.4700 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 309.4550 0.0000 309.5450 0.4700 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 306.8550 0.0000 306.9450 0.4700 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 304.2550 0.0000 304.3450 0.4700 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 301.6550 0.0000 301.7450 0.4700 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 299.0550 0.0000 299.1450 0.4700 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 296.4550 0.0000 296.5450 0.4700 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 293.8550 0.0000 293.9450 0.4700 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 291.2550 0.0000 291.3450 0.4700 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 288.6550 0.0000 288.7450 0.4700 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 286.0550 0.0000 286.1450 0.4700 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 283.4550 0.0000 283.5450 0.4700 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 280.8550 0.0000 280.9450 0.4700 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 278.2550 0.0000 278.3450 0.4700 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 275.6550 0.0000 275.7450 0.4700 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 273.0550 0.0000 273.1450 0.4700 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 270.4550 0.0000 270.5450 0.4700 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 267.8550 0.0000 267.9450 0.4700 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 265.2550 0.0000 265.3450 0.4700 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 262.6550 0.0000 262.7450 0.4700 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 260.0550 0.0000 260.1450 0.4700 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 257.4550 0.0000 257.5450 0.4700 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 254.8550 0.0000 254.9450 0.4700 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 252.2550 0.0000 252.3450 0.4700 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 249.6550 0.0000 249.7450 0.4700 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 247.0550 0.0000 247.1450 0.4700 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 244.4550 0.0000 244.5450 0.4700 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 241.8550 0.0000 241.9450 0.4700 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 239.2550 0.0000 239.3450 0.4700 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 236.6550 0.0000 236.7450 0.4700 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 234.0550 0.0000 234.1450 0.4700 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 231.4550 0.0000 231.5450 0.4700 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 228.8550 0.0000 228.9450 0.4700 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 226.2550 0.0000 226.3450 0.4700 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 223.6550 0.0000 223.7450 0.4700 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 221.0550 0.0000 221.1450 0.4700 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 218.4550 0.0000 218.5450 0.4700 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 215.8550 0.0000 215.9450 0.4700 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 213.2550 0.0000 213.3450 0.4700 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 210.6550 0.0000 210.7450 0.4700 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 208.0550 0.0000 208.1450 0.4700 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 205.4550 0.0000 205.5450 0.4700 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 202.8550 0.0000 202.9450 0.4700 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 200.2550 0.0000 200.3450 0.4700 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 197.6550 0.0000 197.7450 0.4700 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 195.0550 0.0000 195.1450 0.4700 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 192.4550 0.0000 192.5450 0.4700 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 189.8550 0.0000 189.9450 0.4700 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 187.2550 0.0000 187.3450 0.4700 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 184.6550 0.0000 184.7450 0.4700 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 182.0550 0.0000 182.1450 0.4700 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 179.4550 0.0000 179.5450 0.4700 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 176.8550 0.0000 176.9450 0.4700 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 174.2550 0.0000 174.3450 0.4700 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 171.6550 0.0000 171.7450 0.4700 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 169.0550 0.0000 169.1450 0.4700 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 166.4550 0.0000 166.5450 0.4700 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 163.8550 0.0000 163.9450 0.4700 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 161.2550 0.0000 161.3450 0.4700 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 158.6550 0.0000 158.7450 0.4700 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 156.0550 0.0000 156.1450 0.4700 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 153.4550 0.0000 153.5450 0.4700 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 150.8550 0.0000 150.9450 0.4700 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 148.2550 0.0000 148.3450 0.4700 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 145.6550 0.0000 145.7450 0.4700 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 143.0550 0.0000 143.1450 0.4700 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 140.4550 0.0000 140.5450 0.4700 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 137.8550 0.0000 137.9450 0.4700 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 135.2550 0.0000 135.3450 0.4700 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 132.6550 0.0000 132.7450 0.4700 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 130.0550 0.0000 130.1450 0.4700 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 127.4550 0.0000 127.5450 0.4700 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 124.8550 0.0000 124.9450 0.4700 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 122.2550 0.0000 122.3450 0.4700 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 119.6550 0.0000 119.7450 0.4700 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 117.0550 0.0000 117.1450 0.4700 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 114.4550 0.0000 114.5450 0.4700 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 111.8550 0.0000 111.9450 0.4700 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 109.2550 0.0000 109.3450 0.4700 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 106.6550 0.0000 106.7450 0.4700 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 104.0550 0.0000 104.1450 0.4700 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 101.4550 0.0000 101.5450 0.4700 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 98.8550 0.0000 98.9450 0.4700 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 96.2550 0.0000 96.3450 0.4700 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 93.6550 0.0000 93.7450 0.4700 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 91.0550 0.0000 91.1450 0.4700 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 88.4550 0.0000 88.5450 0.4700 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 85.8550 0.0000 85.9450 0.4700 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 83.2550 0.0000 83.3450 0.4700 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 80.6550 0.0000 80.7450 0.4700 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 78.0550 0.0000 78.1450 0.4700 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 122.9500 0.5200 123.0500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 119.9500 0.5200 120.0500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 116.9500 0.5200 117.0500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 113.9500 0.5200 114.0500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 110.9500 0.5200 111.0500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 107.9500 0.5200 108.0500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 104.9500 0.5200 105.0500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 101.9500 0.5200 102.0500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 98.9500 0.5200 99.0500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 95.9500 0.5200 96.0500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 92.9500 0.5200 93.0500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 89.9500 0.5200 90.0500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 86.9500 0.5200 87.0500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 83.9500 0.5200 84.0500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 80.9500 0.5200 81.0500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 77.9500 0.5200 78.0500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 74.9500 0.5200 75.0500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 569.4800 235.1500 570.0000 235.2500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 285.1050 469.3700 570.0000 470.0000 ;
      RECT 0.0000 469.3700 284.6950 470.0000 ;
      RECT 0.0000 0.6300 570.0000 469.3700 ;
      RECT 491.7050 0.0000 570.0000 0.6300 ;
      RECT 489.1050 0.0000 491.2950 0.6300 ;
      RECT 486.5050 0.0000 488.6950 0.6300 ;
      RECT 483.9050 0.0000 486.0950 0.6300 ;
      RECT 481.3050 0.0000 483.4950 0.6300 ;
      RECT 478.7050 0.0000 480.8950 0.6300 ;
      RECT 476.1050 0.0000 478.2950 0.6300 ;
      RECT 473.5050 0.0000 475.6950 0.6300 ;
      RECT 470.9050 0.0000 473.0950 0.6300 ;
      RECT 468.3050 0.0000 470.4950 0.6300 ;
      RECT 465.7050 0.0000 467.8950 0.6300 ;
      RECT 463.1050 0.0000 465.2950 0.6300 ;
      RECT 460.5050 0.0000 462.6950 0.6300 ;
      RECT 457.9050 0.0000 460.0950 0.6300 ;
      RECT 455.3050 0.0000 457.4950 0.6300 ;
      RECT 452.7050 0.0000 454.8950 0.6300 ;
      RECT 450.1050 0.0000 452.2950 0.6300 ;
      RECT 447.5050 0.0000 449.6950 0.6300 ;
      RECT 444.9050 0.0000 447.0950 0.6300 ;
      RECT 442.3050 0.0000 444.4950 0.6300 ;
      RECT 439.7050 0.0000 441.8950 0.6300 ;
      RECT 437.1050 0.0000 439.2950 0.6300 ;
      RECT 434.5050 0.0000 436.6950 0.6300 ;
      RECT 431.9050 0.0000 434.0950 0.6300 ;
      RECT 429.3050 0.0000 431.4950 0.6300 ;
      RECT 426.7050 0.0000 428.8950 0.6300 ;
      RECT 424.1050 0.0000 426.2950 0.6300 ;
      RECT 421.5050 0.0000 423.6950 0.6300 ;
      RECT 418.9050 0.0000 421.0950 0.6300 ;
      RECT 416.3050 0.0000 418.4950 0.6300 ;
      RECT 413.7050 0.0000 415.8950 0.6300 ;
      RECT 411.1050 0.0000 413.2950 0.6300 ;
      RECT 408.5050 0.0000 410.6950 0.6300 ;
      RECT 405.9050 0.0000 408.0950 0.6300 ;
      RECT 403.3050 0.0000 405.4950 0.6300 ;
      RECT 400.7050 0.0000 402.8950 0.6300 ;
      RECT 398.1050 0.0000 400.2950 0.6300 ;
      RECT 395.5050 0.0000 397.6950 0.6300 ;
      RECT 392.9050 0.0000 395.0950 0.6300 ;
      RECT 390.3050 0.0000 392.4950 0.6300 ;
      RECT 387.7050 0.0000 389.8950 0.6300 ;
      RECT 385.1050 0.0000 387.2950 0.6300 ;
      RECT 382.5050 0.0000 384.6950 0.6300 ;
      RECT 379.9050 0.0000 382.0950 0.6300 ;
      RECT 377.3050 0.0000 379.4950 0.6300 ;
      RECT 374.7050 0.0000 376.8950 0.6300 ;
      RECT 372.1050 0.0000 374.2950 0.6300 ;
      RECT 369.5050 0.0000 371.6950 0.6300 ;
      RECT 366.9050 0.0000 369.0950 0.6300 ;
      RECT 364.3050 0.0000 366.4950 0.6300 ;
      RECT 361.7050 0.0000 363.8950 0.6300 ;
      RECT 359.1050 0.0000 361.2950 0.6300 ;
      RECT 356.5050 0.0000 358.6950 0.6300 ;
      RECT 353.9050 0.0000 356.0950 0.6300 ;
      RECT 351.3050 0.0000 353.4950 0.6300 ;
      RECT 348.7050 0.0000 350.8950 0.6300 ;
      RECT 346.1050 0.0000 348.2950 0.6300 ;
      RECT 343.5050 0.0000 345.6950 0.6300 ;
      RECT 340.9050 0.0000 343.0950 0.6300 ;
      RECT 338.3050 0.0000 340.4950 0.6300 ;
      RECT 335.7050 0.0000 337.8950 0.6300 ;
      RECT 333.1050 0.0000 335.2950 0.6300 ;
      RECT 330.5050 0.0000 332.6950 0.6300 ;
      RECT 327.9050 0.0000 330.0950 0.6300 ;
      RECT 325.3050 0.0000 327.4950 0.6300 ;
      RECT 322.7050 0.0000 324.8950 0.6300 ;
      RECT 320.1050 0.0000 322.2950 0.6300 ;
      RECT 317.5050 0.0000 319.6950 0.6300 ;
      RECT 314.9050 0.0000 317.0950 0.6300 ;
      RECT 312.3050 0.0000 314.4950 0.6300 ;
      RECT 309.7050 0.0000 311.8950 0.6300 ;
      RECT 307.1050 0.0000 309.2950 0.6300 ;
      RECT 304.5050 0.0000 306.6950 0.6300 ;
      RECT 301.9050 0.0000 304.0950 0.6300 ;
      RECT 299.3050 0.0000 301.4950 0.6300 ;
      RECT 296.7050 0.0000 298.8950 0.6300 ;
      RECT 294.1050 0.0000 296.2950 0.6300 ;
      RECT 291.5050 0.0000 293.6950 0.6300 ;
      RECT 288.9050 0.0000 291.0950 0.6300 ;
      RECT 286.3050 0.0000 288.4950 0.6300 ;
      RECT 283.7050 0.0000 285.8950 0.6300 ;
      RECT 281.1050 0.0000 283.2950 0.6300 ;
      RECT 278.5050 0.0000 280.6950 0.6300 ;
      RECT 275.9050 0.0000 278.0950 0.6300 ;
      RECT 273.3050 0.0000 275.4950 0.6300 ;
      RECT 270.7050 0.0000 272.8950 0.6300 ;
      RECT 268.1050 0.0000 270.2950 0.6300 ;
      RECT 265.5050 0.0000 267.6950 0.6300 ;
      RECT 262.9050 0.0000 265.0950 0.6300 ;
      RECT 260.3050 0.0000 262.4950 0.6300 ;
      RECT 257.7050 0.0000 259.8950 0.6300 ;
      RECT 255.1050 0.0000 257.2950 0.6300 ;
      RECT 252.5050 0.0000 254.6950 0.6300 ;
      RECT 249.9050 0.0000 252.0950 0.6300 ;
      RECT 247.3050 0.0000 249.4950 0.6300 ;
      RECT 244.7050 0.0000 246.8950 0.6300 ;
      RECT 242.1050 0.0000 244.2950 0.6300 ;
      RECT 239.5050 0.0000 241.6950 0.6300 ;
      RECT 236.9050 0.0000 239.0950 0.6300 ;
      RECT 234.3050 0.0000 236.4950 0.6300 ;
      RECT 231.7050 0.0000 233.8950 0.6300 ;
      RECT 229.1050 0.0000 231.2950 0.6300 ;
      RECT 226.5050 0.0000 228.6950 0.6300 ;
      RECT 223.9050 0.0000 226.0950 0.6300 ;
      RECT 221.3050 0.0000 223.4950 0.6300 ;
      RECT 218.7050 0.0000 220.8950 0.6300 ;
      RECT 216.1050 0.0000 218.2950 0.6300 ;
      RECT 213.5050 0.0000 215.6950 0.6300 ;
      RECT 210.9050 0.0000 213.0950 0.6300 ;
      RECT 208.3050 0.0000 210.4950 0.6300 ;
      RECT 205.7050 0.0000 207.8950 0.6300 ;
      RECT 203.1050 0.0000 205.2950 0.6300 ;
      RECT 200.5050 0.0000 202.6950 0.6300 ;
      RECT 197.9050 0.0000 200.0950 0.6300 ;
      RECT 195.3050 0.0000 197.4950 0.6300 ;
      RECT 192.7050 0.0000 194.8950 0.6300 ;
      RECT 190.1050 0.0000 192.2950 0.6300 ;
      RECT 187.5050 0.0000 189.6950 0.6300 ;
      RECT 184.9050 0.0000 187.0950 0.6300 ;
      RECT 182.3050 0.0000 184.4950 0.6300 ;
      RECT 179.7050 0.0000 181.8950 0.6300 ;
      RECT 177.1050 0.0000 179.2950 0.6300 ;
      RECT 174.5050 0.0000 176.6950 0.6300 ;
      RECT 171.9050 0.0000 174.0950 0.6300 ;
      RECT 169.3050 0.0000 171.4950 0.6300 ;
      RECT 166.7050 0.0000 168.8950 0.6300 ;
      RECT 164.1050 0.0000 166.2950 0.6300 ;
      RECT 161.5050 0.0000 163.6950 0.6300 ;
      RECT 158.9050 0.0000 161.0950 0.6300 ;
      RECT 156.3050 0.0000 158.4950 0.6300 ;
      RECT 153.7050 0.0000 155.8950 0.6300 ;
      RECT 151.1050 0.0000 153.2950 0.6300 ;
      RECT 148.5050 0.0000 150.6950 0.6300 ;
      RECT 145.9050 0.0000 148.0950 0.6300 ;
      RECT 143.3050 0.0000 145.4950 0.6300 ;
      RECT 140.7050 0.0000 142.8950 0.6300 ;
      RECT 138.1050 0.0000 140.2950 0.6300 ;
      RECT 135.5050 0.0000 137.6950 0.6300 ;
      RECT 132.9050 0.0000 135.0950 0.6300 ;
      RECT 130.3050 0.0000 132.4950 0.6300 ;
      RECT 127.7050 0.0000 129.8950 0.6300 ;
      RECT 125.1050 0.0000 127.2950 0.6300 ;
      RECT 122.5050 0.0000 124.6950 0.6300 ;
      RECT 119.9050 0.0000 122.0950 0.6300 ;
      RECT 117.3050 0.0000 119.4950 0.6300 ;
      RECT 114.7050 0.0000 116.8950 0.6300 ;
      RECT 112.1050 0.0000 114.2950 0.6300 ;
      RECT 109.5050 0.0000 111.6950 0.6300 ;
      RECT 106.9050 0.0000 109.0950 0.6300 ;
      RECT 104.3050 0.0000 106.4950 0.6300 ;
      RECT 101.7050 0.0000 103.8950 0.6300 ;
      RECT 99.1050 0.0000 101.2950 0.6300 ;
      RECT 96.5050 0.0000 98.6950 0.6300 ;
      RECT 93.9050 0.0000 96.0950 0.6300 ;
      RECT 91.3050 0.0000 93.4950 0.6300 ;
      RECT 88.7050 0.0000 90.8950 0.6300 ;
      RECT 86.1050 0.0000 88.2950 0.6300 ;
      RECT 83.5050 0.0000 85.6950 0.6300 ;
      RECT 80.9050 0.0000 83.0950 0.6300 ;
      RECT 78.3050 0.0000 80.4950 0.6300 ;
      RECT 0.0000 0.0000 77.8950 0.6300 ;
    LAYER M2 ;
      RECT 0.0000 315.2100 570.0000 470.0000 ;
      RECT 0.6800 314.7900 570.0000 315.2100 ;
      RECT 0.0000 312.2100 570.0000 314.7900 ;
      RECT 0.6800 311.7900 570.0000 312.2100 ;
      RECT 0.0000 309.2100 570.0000 311.7900 ;
      RECT 0.6800 308.7900 570.0000 309.2100 ;
      RECT 0.0000 306.2100 570.0000 308.7900 ;
      RECT 0.6800 305.7900 570.0000 306.2100 ;
      RECT 0.0000 303.2100 570.0000 305.7900 ;
      RECT 0.6800 302.7900 570.0000 303.2100 ;
      RECT 0.0000 300.2100 570.0000 302.7900 ;
      RECT 0.6800 299.7900 570.0000 300.2100 ;
      RECT 0.0000 297.2100 570.0000 299.7900 ;
      RECT 0.6800 296.7900 570.0000 297.2100 ;
      RECT 0.0000 294.2100 570.0000 296.7900 ;
      RECT 0.6800 293.7900 570.0000 294.2100 ;
      RECT 0.0000 291.2100 570.0000 293.7900 ;
      RECT 0.6800 290.7900 570.0000 291.2100 ;
      RECT 0.0000 288.2100 570.0000 290.7900 ;
      RECT 0.6800 287.7900 570.0000 288.2100 ;
      RECT 0.0000 285.2100 570.0000 287.7900 ;
      RECT 0.6800 284.7900 570.0000 285.2100 ;
      RECT 0.0000 282.2100 570.0000 284.7900 ;
      RECT 0.6800 281.7900 570.0000 282.2100 ;
      RECT 0.0000 279.2100 570.0000 281.7900 ;
      RECT 0.6800 278.7900 570.0000 279.2100 ;
      RECT 0.0000 276.2100 570.0000 278.7900 ;
      RECT 0.6800 275.7900 570.0000 276.2100 ;
      RECT 0.0000 273.2100 570.0000 275.7900 ;
      RECT 0.6800 272.7900 570.0000 273.2100 ;
      RECT 0.0000 270.2100 570.0000 272.7900 ;
      RECT 0.6800 269.7900 570.0000 270.2100 ;
      RECT 0.0000 267.2100 570.0000 269.7900 ;
      RECT 0.6800 266.7900 570.0000 267.2100 ;
      RECT 0.0000 264.2100 570.0000 266.7900 ;
      RECT 0.6800 263.7900 570.0000 264.2100 ;
      RECT 0.0000 261.2100 570.0000 263.7900 ;
      RECT 0.6800 260.7900 570.0000 261.2100 ;
      RECT 0.0000 258.2100 570.0000 260.7900 ;
      RECT 0.6800 257.7900 570.0000 258.2100 ;
      RECT 0.0000 255.2100 570.0000 257.7900 ;
      RECT 0.6800 254.7900 570.0000 255.2100 ;
      RECT 0.0000 252.2100 570.0000 254.7900 ;
      RECT 0.6800 251.7900 570.0000 252.2100 ;
      RECT 0.0000 249.2100 570.0000 251.7900 ;
      RECT 0.6800 248.7900 570.0000 249.2100 ;
      RECT 0.0000 246.2100 570.0000 248.7900 ;
      RECT 0.6800 245.7900 570.0000 246.2100 ;
      RECT 0.0000 243.2100 570.0000 245.7900 ;
      RECT 0.6800 242.7900 570.0000 243.2100 ;
      RECT 0.0000 240.2100 570.0000 242.7900 ;
      RECT 0.6800 239.7900 570.0000 240.2100 ;
      RECT 0.0000 237.2100 570.0000 239.7900 ;
      RECT 0.6800 236.7900 570.0000 237.2100 ;
      RECT 0.0000 235.4100 570.0000 236.7900 ;
      RECT 0.0000 234.9900 569.3200 235.4100 ;
      RECT 0.0000 234.2100 570.0000 234.9900 ;
      RECT 0.6800 233.7900 570.0000 234.2100 ;
      RECT 0.0000 231.2100 570.0000 233.7900 ;
      RECT 0.6800 230.7900 570.0000 231.2100 ;
      RECT 0.0000 228.2100 570.0000 230.7900 ;
      RECT 0.6800 227.7900 570.0000 228.2100 ;
      RECT 0.0000 225.2100 570.0000 227.7900 ;
      RECT 0.6800 224.7900 570.0000 225.2100 ;
      RECT 0.0000 222.2100 570.0000 224.7900 ;
      RECT 0.6800 221.7900 570.0000 222.2100 ;
      RECT 0.0000 219.2100 570.0000 221.7900 ;
      RECT 0.6800 218.7900 570.0000 219.2100 ;
      RECT 0.0000 216.2100 570.0000 218.7900 ;
      RECT 0.6800 215.7900 570.0000 216.2100 ;
      RECT 0.0000 213.2100 570.0000 215.7900 ;
      RECT 0.6800 212.7900 570.0000 213.2100 ;
      RECT 0.0000 210.2100 570.0000 212.7900 ;
      RECT 0.6800 209.7900 570.0000 210.2100 ;
      RECT 0.0000 207.2100 570.0000 209.7900 ;
      RECT 0.6800 206.7900 570.0000 207.2100 ;
      RECT 0.0000 204.2100 570.0000 206.7900 ;
      RECT 0.6800 203.7900 570.0000 204.2100 ;
      RECT 0.0000 201.2100 570.0000 203.7900 ;
      RECT 0.6800 200.7900 570.0000 201.2100 ;
      RECT 0.0000 198.2100 570.0000 200.7900 ;
      RECT 0.6800 197.7900 570.0000 198.2100 ;
      RECT 0.0000 195.2100 570.0000 197.7900 ;
      RECT 0.6800 194.7900 570.0000 195.2100 ;
      RECT 0.0000 192.2100 570.0000 194.7900 ;
      RECT 0.6800 191.7900 570.0000 192.2100 ;
      RECT 0.0000 189.2100 570.0000 191.7900 ;
      RECT 0.6800 188.7900 570.0000 189.2100 ;
      RECT 0.0000 186.2100 570.0000 188.7900 ;
      RECT 0.6800 185.7900 570.0000 186.2100 ;
      RECT 0.0000 183.2100 570.0000 185.7900 ;
      RECT 0.6800 182.7900 570.0000 183.2100 ;
      RECT 0.0000 180.2100 570.0000 182.7900 ;
      RECT 0.6800 179.7900 570.0000 180.2100 ;
      RECT 0.0000 177.2100 570.0000 179.7900 ;
      RECT 0.6800 176.7900 570.0000 177.2100 ;
      RECT 0.0000 174.2100 570.0000 176.7900 ;
      RECT 0.6800 173.7900 570.0000 174.2100 ;
      RECT 0.0000 171.2100 570.0000 173.7900 ;
      RECT 0.6800 170.7900 570.0000 171.2100 ;
      RECT 0.0000 168.2100 570.0000 170.7900 ;
      RECT 0.6800 167.7900 570.0000 168.2100 ;
      RECT 0.0000 165.2100 570.0000 167.7900 ;
      RECT 0.6800 164.7900 570.0000 165.2100 ;
      RECT 0.0000 162.2100 570.0000 164.7900 ;
      RECT 0.6800 161.7900 570.0000 162.2100 ;
      RECT 0.0000 159.2100 570.0000 161.7900 ;
      RECT 0.6800 158.7900 570.0000 159.2100 ;
      RECT 0.0000 156.2100 570.0000 158.7900 ;
      RECT 0.6800 155.7900 570.0000 156.2100 ;
      RECT 0.0000 153.2100 570.0000 155.7900 ;
      RECT 0.6800 152.7900 570.0000 153.2100 ;
      RECT 0.0000 150.2100 570.0000 152.7900 ;
      RECT 0.6800 149.7900 570.0000 150.2100 ;
      RECT 0.0000 147.2100 570.0000 149.7900 ;
      RECT 0.6800 146.7900 570.0000 147.2100 ;
      RECT 0.0000 144.2100 570.0000 146.7900 ;
      RECT 0.6800 143.7900 570.0000 144.2100 ;
      RECT 0.0000 141.2100 570.0000 143.7900 ;
      RECT 0.6800 140.7900 570.0000 141.2100 ;
      RECT 0.0000 138.2100 570.0000 140.7900 ;
      RECT 0.6800 137.7900 570.0000 138.2100 ;
      RECT 0.0000 135.2100 570.0000 137.7900 ;
      RECT 0.6800 134.7900 570.0000 135.2100 ;
      RECT 0.0000 132.2100 570.0000 134.7900 ;
      RECT 0.6800 131.7900 570.0000 132.2100 ;
      RECT 0.0000 129.2100 570.0000 131.7900 ;
      RECT 0.6800 128.7900 570.0000 129.2100 ;
      RECT 0.0000 126.2100 570.0000 128.7900 ;
      RECT 0.6800 125.7900 570.0000 126.2100 ;
      RECT 0.0000 123.2100 570.0000 125.7900 ;
      RECT 0.6800 122.7900 570.0000 123.2100 ;
      RECT 0.0000 120.2100 570.0000 122.7900 ;
      RECT 0.6800 119.7900 570.0000 120.2100 ;
      RECT 0.0000 117.2100 570.0000 119.7900 ;
      RECT 0.6800 116.7900 570.0000 117.2100 ;
      RECT 0.0000 114.2100 570.0000 116.7900 ;
      RECT 0.6800 113.7900 570.0000 114.2100 ;
      RECT 0.0000 111.2100 570.0000 113.7900 ;
      RECT 0.6800 110.7900 570.0000 111.2100 ;
      RECT 0.0000 108.2100 570.0000 110.7900 ;
      RECT 0.6800 107.7900 570.0000 108.2100 ;
      RECT 0.0000 105.2100 570.0000 107.7900 ;
      RECT 0.6800 104.7900 570.0000 105.2100 ;
      RECT 0.0000 102.2100 570.0000 104.7900 ;
      RECT 0.6800 101.7900 570.0000 102.2100 ;
      RECT 0.0000 99.2100 570.0000 101.7900 ;
      RECT 0.6800 98.7900 570.0000 99.2100 ;
      RECT 0.0000 96.2100 570.0000 98.7900 ;
      RECT 0.6800 95.7900 570.0000 96.2100 ;
      RECT 0.0000 93.2100 570.0000 95.7900 ;
      RECT 0.6800 92.7900 570.0000 93.2100 ;
      RECT 0.0000 90.2100 570.0000 92.7900 ;
      RECT 0.6800 89.7900 570.0000 90.2100 ;
      RECT 0.0000 87.2100 570.0000 89.7900 ;
      RECT 0.6800 86.7900 570.0000 87.2100 ;
      RECT 0.0000 84.2100 570.0000 86.7900 ;
      RECT 0.6800 83.7900 570.0000 84.2100 ;
      RECT 0.0000 81.2100 570.0000 83.7900 ;
      RECT 0.6800 80.7900 570.0000 81.2100 ;
      RECT 0.0000 78.2100 570.0000 80.7900 ;
      RECT 0.6800 77.7900 570.0000 78.2100 ;
      RECT 0.0000 75.2100 570.0000 77.7900 ;
      RECT 0.6800 74.7900 570.0000 75.2100 ;
      RECT 0.0000 0.0000 570.0000 74.7900 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 570.0000 470.0000 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 570.0000 470.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 570.0000 470.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 570.0000 470.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 570.0000 470.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 570.0000 470.0000 ;
  END
END core

END LIBRARY
