##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Wed Mar 19 22:02:05 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 1120.0000 BY 1120.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.8500 1119.4800 395.9500 1120.0000 ;
    END
  END clk
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.0500 0.0000 194.1500 0.5200 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.0500 0.0000 198.1500 0.5200 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.0500 0.0000 202.1500 0.5200 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.0500 0.0000 206.1500 0.5200 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.0500 0.0000 210.1500 0.5200 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.0500 0.0000 214.1500 0.5200 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.0500 0.0000 218.1500 0.5200 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.0500 0.0000 222.1500 0.5200 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.0500 0.0000 226.1500 0.5200 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.0500 0.0000 230.1500 0.5200 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.0500 0.0000 234.1500 0.5200 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.0500 0.0000 238.1500 0.5200 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 242.0500 0.0000 242.1500 0.5200 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.0500 0.0000 246.1500 0.5200 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.0500 0.0000 250.1500 0.5200 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 254.0500 0.0000 254.1500 0.5200 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.0500 0.0000 258.1500 0.5200 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.0500 0.0000 262.1500 0.5200 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 266.0500 0.0000 266.1500 0.5200 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.0500 0.0000 270.1500 0.5200 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.0500 0.0000 274.1500 0.5200 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.0500 0.0000 278.1500 0.5200 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.0500 0.0000 282.1500 0.5200 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 286.0500 0.0000 286.1500 0.5200 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 719.8500 1119.4800 719.9500 1120.0000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 715.8500 1119.4800 715.9500 1120.0000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 711.8500 1119.4800 711.9500 1120.0000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 707.8500 1119.4800 707.9500 1120.0000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 703.8500 1119.4800 703.9500 1120.0000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 699.8500 1119.4800 699.9500 1120.0000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 695.8500 1119.4800 695.9500 1120.0000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 691.8500 1119.4800 691.9500 1120.0000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 687.8500 1119.4800 687.9500 1120.0000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 683.8500 1119.4800 683.9500 1120.0000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 679.8500 1119.4800 679.9500 1120.0000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 675.8500 1119.4800 675.9500 1120.0000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 671.8500 1119.4800 671.9500 1120.0000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 667.8500 1119.4800 667.9500 1120.0000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 663.8500 1119.4800 663.9500 1120.0000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 659.8500 1119.4800 659.9500 1120.0000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 655.8500 1119.4800 655.9500 1120.0000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 651.8500 1119.4800 651.9500 1120.0000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 647.8500 1119.4800 647.9500 1120.0000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 643.8500 1119.4800 643.9500 1120.0000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 639.8500 1119.4800 639.9500 1120.0000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 635.8500 1119.4800 635.9500 1120.0000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 631.8500 1119.4800 631.9500 1120.0000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 627.8500 1119.4800 627.9500 1120.0000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 623.8500 1119.4800 623.9500 1120.0000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 619.8500 1119.4800 619.9500 1120.0000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 615.8500 1119.4800 615.9500 1120.0000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 611.8500 1119.4800 611.9500 1120.0000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 607.8500 1119.4800 607.9500 1120.0000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 603.8500 1119.4800 603.9500 1120.0000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 599.8500 1119.4800 599.9500 1120.0000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 595.8500 1119.4800 595.9500 1120.0000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 591.8500 1119.4800 591.9500 1120.0000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 587.8500 1119.4800 587.9500 1120.0000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 583.8500 1119.4800 583.9500 1120.0000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 579.8500 1119.4800 579.9500 1120.0000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 575.8500 1119.4800 575.9500 1120.0000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 571.8500 1119.4800 571.9500 1120.0000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 567.8500 1119.4800 567.9500 1120.0000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 563.8500 1119.4800 563.9500 1120.0000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 559.8500 1119.4800 559.9500 1120.0000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 555.8500 1119.4800 555.9500 1120.0000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 551.8500 1119.4800 551.9500 1120.0000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 547.8500 1119.4800 547.9500 1120.0000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 543.8500 1119.4800 543.9500 1120.0000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 539.8500 1119.4800 539.9500 1120.0000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 535.8500 1119.4800 535.9500 1120.0000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 531.8500 1119.4800 531.9500 1120.0000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 527.8500 1119.4800 527.9500 1120.0000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 523.8500 1119.4800 523.9500 1120.0000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 519.8500 1119.4800 519.9500 1120.0000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 515.8500 1119.4800 515.9500 1120.0000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 511.8500 1119.4800 511.9500 1120.0000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.8500 1119.4800 507.9500 1120.0000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 503.8500 1119.4800 503.9500 1120.0000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 499.8500 1119.4800 499.9500 1120.0000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 495.8500 1119.4800 495.9500 1120.0000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 491.8500 1119.4800 491.9500 1120.0000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 487.8500 1119.4800 487.9500 1120.0000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 483.8500 1119.4800 483.9500 1120.0000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 479.8500 1119.4800 479.9500 1120.0000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 475.8500 1119.4800 475.9500 1120.0000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 471.8500 1119.4800 471.9500 1120.0000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 467.8500 1119.4800 467.9500 1120.0000 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 290.0500 0.0000 290.1500 0.5200 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 294.0500 0.0000 294.1500 0.5200 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 298.0500 0.0000 298.1500 0.5200 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.0500 0.0000 302.1500 0.5200 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.0500 0.0000 306.1500 0.5200 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.0500 0.0000 310.1500 0.5200 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.0500 0.0000 314.1500 0.5200 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.0500 0.0000 318.1500 0.5200 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.0500 0.0000 322.1500 0.5200 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.0500 0.0000 326.1500 0.5200 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.0500 0.0000 330.1500 0.5200 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.0500 0.0000 334.1500 0.5200 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.0500 0.0000 338.1500 0.5200 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.0500 0.0000 342.1500 0.5200 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.0500 0.0000 346.1500 0.5200 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.0500 0.0000 350.1500 0.5200 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.0500 0.0000 354.1500 0.5200 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.0500 0.0000 358.1500 0.5200 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.0500 0.0000 362.1500 0.5200 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.0500 0.0000 366.1500 0.5200 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.0500 0.0000 370.1500 0.5200 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.0500 0.0000 374.1500 0.5200 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.0500 0.0000 378.1500 0.5200 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.0500 0.0000 382.1500 0.5200 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.0500 0.0000 386.1500 0.5200 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.0500 0.0000 390.1500 0.5200 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.0500 0.0000 394.1500 0.5200 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.0500 0.0000 398.1500 0.5200 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.0500 0.0000 402.1500 0.5200 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.0500 0.0000 406.1500 0.5200 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.0500 0.0000 410.1500 0.5200 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.0500 0.0000 414.1500 0.5200 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.0500 0.0000 418.1500 0.5200 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.0500 0.0000 422.1500 0.5200 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.0500 0.0000 426.1500 0.5200 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.0500 0.0000 430.1500 0.5200 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.0500 0.0000 434.1500 0.5200 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.0500 0.0000 438.1500 0.5200 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.0500 0.0000 442.1500 0.5200 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.0500 0.0000 446.1500 0.5200 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.0500 0.0000 450.1500 0.5200 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.0500 0.0000 454.1500 0.5200 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 458.0500 0.0000 458.1500 0.5200 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 462.0500 0.0000 462.1500 0.5200 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 466.0500 0.0000 466.1500 0.5200 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 470.0500 0.0000 470.1500 0.5200 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 474.0500 0.0000 474.1500 0.5200 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 478.0500 0.0000 478.1500 0.5200 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 482.0500 0.0000 482.1500 0.5200 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 486.0500 0.0000 486.1500 0.5200 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 490.0500 0.0000 490.1500 0.5200 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 494.0500 0.0000 494.1500 0.5200 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 498.0500 0.0000 498.1500 0.5200 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 502.0500 0.0000 502.1500 0.5200 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 506.0500 0.0000 506.1500 0.5200 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 510.0500 0.0000 510.1500 0.5200 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 514.0500 0.0000 514.1500 0.5200 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 518.0500 0.0000 518.1500 0.5200 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 522.0500 0.0000 522.1500 0.5200 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 526.0500 0.0000 526.1500 0.5200 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 530.0500 0.0000 530.1500 0.5200 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 534.0500 0.0000 534.1500 0.5200 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 538.0500 0.0000 538.1500 0.5200 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 542.0500 0.0000 542.1500 0.5200 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 546.0500 0.0000 546.1500 0.5200 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 550.0500 0.0000 550.1500 0.5200 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 554.0500 0.0000 554.1500 0.5200 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 558.0500 0.0000 558.1500 0.5200 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 562.0500 0.0000 562.1500 0.5200 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 566.0500 0.0000 566.1500 0.5200 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 570.0500 0.0000 570.1500 0.5200 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 574.0500 0.0000 574.1500 0.5200 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 578.0500 0.0000 578.1500 0.5200 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 582.0500 0.0000 582.1500 0.5200 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 586.0500 0.0000 586.1500 0.5200 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 590.0500 0.0000 590.1500 0.5200 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 594.0500 0.0000 594.1500 0.5200 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 598.0500 0.0000 598.1500 0.5200 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 602.0500 0.0000 602.1500 0.5200 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 606.0500 0.0000 606.1500 0.5200 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 610.0500 0.0000 610.1500 0.5200 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 614.0500 0.0000 614.1500 0.5200 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 618.0500 0.0000 618.1500 0.5200 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 622.0500 0.0000 622.1500 0.5200 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 626.0500 0.0000 626.1500 0.5200 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 630.0500 0.0000 630.1500 0.5200 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 634.0500 0.0000 634.1500 0.5200 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 638.0500 0.0000 638.1500 0.5200 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 642.0500 0.0000 642.1500 0.5200 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 646.0500 0.0000 646.1500 0.5200 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 650.0500 0.0000 650.1500 0.5200 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 654.0500 0.0000 654.1500 0.5200 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 658.0500 0.0000 658.1500 0.5200 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 662.0500 0.0000 662.1500 0.5200 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 666.0500 0.0000 666.1500 0.5200 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 670.0500 0.0000 670.1500 0.5200 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 674.0500 0.0000 674.1500 0.5200 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 678.0500 0.0000 678.1500 0.5200 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 682.0500 0.0000 682.1500 0.5200 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 686.0500 0.0000 686.1500 0.5200 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690.0500 0.0000 690.1500 0.5200 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 694.0500 0.0000 694.1500 0.5200 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 698.0500 0.0000 698.1500 0.5200 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 702.0500 0.0000 702.1500 0.5200 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 706.0500 0.0000 706.1500 0.5200 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 710.0500 0.0000 710.1500 0.5200 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 714.0500 0.0000 714.1500 0.5200 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 718.0500 0.0000 718.1500 0.5200 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 722.0500 0.0000 722.1500 0.5200 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 726.0500 0.0000 726.1500 0.5200 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 730.0500 0.0000 730.1500 0.5200 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 734.0500 0.0000 734.1500 0.5200 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 738.0500 0.0000 738.1500 0.5200 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 742.0500 0.0000 742.1500 0.5200 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 746.0500 0.0000 746.1500 0.5200 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 750.0500 0.0000 750.1500 0.5200 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 754.0500 0.0000 754.1500 0.5200 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 758.0500 0.0000 758.1500 0.5200 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 762.0500 0.0000 762.1500 0.5200 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 766.0500 0.0000 766.1500 0.5200 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 770.0500 0.0000 770.1500 0.5200 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 774.0500 0.0000 774.1500 0.5200 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 778.0500 0.0000 778.1500 0.5200 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 782.0500 0.0000 782.1500 0.5200 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 786.0500 0.0000 786.1500 0.5200 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 790.0500 0.0000 790.1500 0.5200 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 794.0500 0.0000 794.1500 0.5200 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 798.0500 0.0000 798.1500 0.5200 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 802.0500 0.0000 802.1500 0.5200 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 806.0500 0.0000 806.1500 0.5200 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 810.0500 0.0000 810.1500 0.5200 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 814.0500 0.0000 814.1500 0.5200 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 818.0500 0.0000 818.1500 0.5200 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 822.0500 0.0000 822.1500 0.5200 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 826.0500 0.0000 826.1500 0.5200 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 830.0500 0.0000 830.1500 0.5200 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 834.0500 0.0000 834.1500 0.5200 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 838.0500 0.0000 838.1500 0.5200 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 842.0500 0.0000 842.1500 0.5200 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 846.0500 0.0000 846.1500 0.5200 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 850.0500 0.0000 850.1500 0.5200 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 854.0500 0.0000 854.1500 0.5200 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 858.0500 0.0000 858.1500 0.5200 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 862.0500 0.0000 862.1500 0.5200 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 866.0500 0.0000 866.1500 0.5200 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 870.0500 0.0000 870.1500 0.5200 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 874.0500 0.0000 874.1500 0.5200 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 878.0500 0.0000 878.1500 0.5200 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 882.0500 0.0000 882.1500 0.5200 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 886.0500 0.0000 886.1500 0.5200 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 890.0500 0.0000 890.1500 0.5200 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 894.0500 0.0000 894.1500 0.5200 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 898.0500 0.0000 898.1500 0.5200 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 902.0500 0.0000 902.1500 0.5200 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 906.0500 0.0000 906.1500 0.5200 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 910.0500 0.0000 910.1500 0.5200 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 914.0500 0.0000 914.1500 0.5200 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 918.0500 0.0000 918.1500 0.5200 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 922.0500 0.0000 922.1500 0.5200 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 926.0500 0.0000 926.1500 0.5200 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.8500 1119.4800 463.9500 1120.0000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 459.8500 1119.4800 459.9500 1120.0000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.8500 1119.4800 455.9500 1120.0000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.8500 1119.4800 451.9500 1120.0000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.8500 1119.4800 447.9500 1120.0000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.8500 1119.4800 443.9500 1120.0000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.8500 1119.4800 439.9500 1120.0000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.8500 1119.4800 435.9500 1120.0000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.8500 1119.4800 431.9500 1120.0000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.8500 1119.4800 427.9500 1120.0000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.8500 1119.4800 423.9500 1120.0000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.8500 1119.4800 419.9500 1120.0000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.8500 1119.4800 415.9500 1120.0000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.8500 1119.4800 411.9500 1120.0000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.8500 1119.4800 407.9500 1120.0000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.8500 1119.4800 403.9500 1120.0000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.8500 1119.4800 399.9500 1120.0000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 723.8500 1119.4800 723.9500 1120.0000 ;
    END
  END reset
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 68.5150 64.6650 70.5150 66.6650 ;
        RECT 6.0000 15.0000 8.0000 17.0000 ;
        RECT 6.0000 22.0950 8.0000 24.0950 ;
        RECT 6.0000 29.1900 8.0000 31.1900 ;
        RECT 6.0000 43.3800 8.0000 45.3800 ;
        RECT 6.0000 36.2850 8.0000 38.2850 ;
        RECT 6.0000 50.4750 8.0000 52.4750 ;
        RECT 6.0000 57.5700 8.0000 59.5700 ;
        RECT 6.0000 64.6650 8.0000 66.6650 ;
        RECT 44.0000 50.4750 46.0000 52.4750 ;
        RECT 44.0000 44.0000 46.0000 45.3800 ;
        RECT 44.0000 57.5700 46.0000 59.5700 ;
        RECT 44.0000 64.6650 46.0000 66.6650 ;
        RECT 60.0000 64.6650 62.0000 66.6650 ;
        RECT 60.0000 60.0000 62.0000 62.0000 ;
        RECT 77.0300 64.6650 79.0300 66.6650 ;
        RECT 85.5450 64.6650 87.5450 66.6650 ;
        RECT 94.0600 64.6650 96.0600 66.6650 ;
        RECT 102.5750 64.6650 104.5750 66.6650 ;
        RECT 111.0900 64.6650 113.0900 66.6650 ;
        RECT 119.6050 64.6650 121.6050 66.6650 ;
        RECT 128.1200 64.6650 130.1200 66.6650 ;
        RECT 136.6350 64.6650 138.6350 66.6650 ;
        RECT 68.5150 71.7600 70.5150 73.7600 ;
        RECT 68.5150 78.8550 70.5150 80.8550 ;
        RECT 68.5150 85.9500 70.5150 87.9500 ;
        RECT 68.5150 93.0450 70.5150 95.0450 ;
        RECT 68.5150 100.1400 70.5150 102.1400 ;
        RECT 68.5150 107.2350 70.5150 109.2350 ;
        RECT 68.5150 114.3300 70.5150 116.3300 ;
        RECT 68.5150 121.4250 70.5150 123.4250 ;
        RECT 68.5150 128.5200 70.5150 130.5200 ;
        RECT 68.5150 135.6150 70.5150 137.6150 ;
        RECT 6.0000 85.9500 8.0000 87.9500 ;
        RECT 6.0000 78.8550 8.0000 80.8550 ;
        RECT 6.0000 71.7600 8.0000 73.7600 ;
        RECT 6.0000 100.1400 8.0000 102.1400 ;
        RECT 6.0000 93.0450 8.0000 95.0450 ;
        RECT 44.0000 85.9500 46.0000 87.9500 ;
        RECT 60.0000 85.9500 62.0000 87.9500 ;
        RECT 44.0000 78.8550 46.0000 80.8550 ;
        RECT 44.0000 71.7600 46.0000 73.7600 ;
        RECT 60.0000 71.7600 62.0000 73.7600 ;
        RECT 60.0000 78.8550 62.0000 80.8550 ;
        RECT 44.0000 100.1400 46.0000 102.1400 ;
        RECT 44.0000 93.0450 46.0000 95.0450 ;
        RECT 60.0000 93.0450 62.0000 95.0450 ;
        RECT 60.0000 100.1400 62.0000 102.1400 ;
        RECT 6.0000 121.4250 8.0000 123.4250 ;
        RECT 6.0000 107.2350 8.0000 109.2350 ;
        RECT 6.0000 114.3300 8.0000 116.3300 ;
        RECT 6.0000 128.5200 8.0000 130.5200 ;
        RECT 6.0000 135.6150 8.0000 137.6150 ;
        RECT 44.0000 121.4250 46.0000 123.4250 ;
        RECT 60.0000 121.4250 62.0000 123.4250 ;
        RECT 44.0000 107.2350 46.0000 109.2350 ;
        RECT 44.0000 114.3300 46.0000 116.3300 ;
        RECT 60.0000 114.3300 62.0000 116.3300 ;
        RECT 60.0000 107.2350 62.0000 109.2350 ;
        RECT 44.0000 128.5200 46.0000 130.5200 ;
        RECT 44.0000 135.6150 46.0000 137.6150 ;
        RECT 60.0000 135.6150 62.0000 137.6150 ;
        RECT 60.0000 128.5200 62.0000 130.5200 ;
        RECT 77.0300 85.9500 79.0300 87.9500 ;
        RECT 85.5450 85.9500 87.5450 87.9500 ;
        RECT 94.0600 85.9500 96.0600 87.9500 ;
        RECT 102.5750 85.9500 104.5750 87.9500 ;
        RECT 102.5750 78.8550 104.5750 80.8550 ;
        RECT 94.0600 78.8550 96.0600 80.8550 ;
        RECT 85.5450 78.8550 87.5450 80.8550 ;
        RECT 77.0300 78.8550 79.0300 80.8550 ;
        RECT 102.5750 71.7600 104.5750 73.7600 ;
        RECT 94.0600 71.7600 96.0600 73.7600 ;
        RECT 85.5450 71.7600 87.5450 73.7600 ;
        RECT 77.0300 71.7600 79.0300 73.7600 ;
        RECT 77.0300 93.0450 79.0300 95.0450 ;
        RECT 85.5450 93.0450 87.5450 95.0450 ;
        RECT 94.0600 93.0450 96.0600 95.0450 ;
        RECT 102.5750 93.0450 104.5750 95.0450 ;
        RECT 77.0300 100.1400 79.0300 102.1400 ;
        RECT 85.5450 100.1400 87.5450 102.1400 ;
        RECT 94.0600 100.1400 96.0600 102.1400 ;
        RECT 102.5750 100.1400 104.5750 102.1400 ;
        RECT 111.0900 85.9500 113.0900 87.9500 ;
        RECT 119.6050 85.9500 121.6050 87.9500 ;
        RECT 128.1200 85.9500 130.1200 87.9500 ;
        RECT 136.6350 85.9500 138.6350 87.9500 ;
        RECT 136.6350 78.8550 138.6350 80.8550 ;
        RECT 128.1200 78.8550 130.1200 80.8550 ;
        RECT 119.6050 78.8550 121.6050 80.8550 ;
        RECT 111.0900 78.8550 113.0900 80.8550 ;
        RECT 136.6350 71.7600 138.6350 73.7600 ;
        RECT 128.1200 71.7600 130.1200 73.7600 ;
        RECT 119.6050 71.7600 121.6050 73.7600 ;
        RECT 111.0900 71.7600 113.0900 73.7600 ;
        RECT 111.0900 93.0450 113.0900 95.0450 ;
        RECT 119.6050 93.0450 121.6050 95.0450 ;
        RECT 128.1200 93.0450 130.1200 95.0450 ;
        RECT 136.6350 93.0450 138.6350 95.0450 ;
        RECT 111.0900 100.1400 113.0900 102.1400 ;
        RECT 119.6050 100.1400 121.6050 102.1400 ;
        RECT 128.1200 100.1400 130.1200 102.1400 ;
        RECT 136.6350 100.1400 138.6350 102.1400 ;
        RECT 77.0300 121.4250 79.0300 123.4250 ;
        RECT 85.5450 121.4250 87.5450 123.4250 ;
        RECT 94.0600 121.4250 96.0600 123.4250 ;
        RECT 102.5750 121.4250 104.5750 123.4250 ;
        RECT 102.5750 114.3300 104.5750 116.3300 ;
        RECT 94.0600 114.3300 96.0600 116.3300 ;
        RECT 85.5450 114.3300 87.5450 116.3300 ;
        RECT 77.0300 114.3300 79.0300 116.3300 ;
        RECT 102.5750 107.2350 104.5750 109.2350 ;
        RECT 94.0600 107.2350 96.0600 109.2350 ;
        RECT 85.5450 107.2350 87.5450 109.2350 ;
        RECT 77.0300 107.2350 79.0300 109.2350 ;
        RECT 77.0300 128.5200 79.0300 130.5200 ;
        RECT 85.5450 128.5200 87.5450 130.5200 ;
        RECT 94.0600 128.5200 96.0600 130.5200 ;
        RECT 102.5750 128.5200 104.5750 130.5200 ;
        RECT 77.0300 135.6150 79.0300 137.6150 ;
        RECT 85.5450 135.6150 87.5450 137.6150 ;
        RECT 94.0600 135.6150 96.0600 137.6150 ;
        RECT 102.5750 135.6150 104.5750 137.6150 ;
        RECT 111.0900 121.4250 113.0900 123.4250 ;
        RECT 119.6050 121.4250 121.6050 123.4250 ;
        RECT 128.1200 121.4250 130.1200 123.4250 ;
        RECT 136.6350 121.4250 138.6350 123.4250 ;
        RECT 136.6350 114.3300 138.6350 116.3300 ;
        RECT 128.1200 114.3300 130.1200 116.3300 ;
        RECT 119.6050 114.3300 121.6050 116.3300 ;
        RECT 111.0900 114.3300 113.0900 116.3300 ;
        RECT 136.6350 107.2350 138.6350 109.2350 ;
        RECT 128.1200 107.2350 130.1200 109.2350 ;
        RECT 119.6050 107.2350 121.6050 109.2350 ;
        RECT 111.0900 107.2350 113.0900 109.2350 ;
        RECT 111.0900 128.5200 113.0900 130.5200 ;
        RECT 119.6050 128.5200 121.6050 130.5200 ;
        RECT 128.1200 128.5200 130.1200 130.5200 ;
        RECT 136.6350 128.5200 138.6350 130.5200 ;
        RECT 111.0900 135.6150 113.0900 137.6150 ;
        RECT 119.6050 135.6150 121.6050 137.6150 ;
        RECT 128.1200 135.6150 130.1200 137.6150 ;
        RECT 136.6350 135.6150 138.6350 137.6150 ;
        RECT 204.7550 64.6650 206.7550 66.6650 ;
        RECT 196.2400 64.6650 198.2400 66.6650 ;
        RECT 187.7250 64.6650 189.7250 66.6650 ;
        RECT 179.2100 64.6650 181.2100 66.6650 ;
        RECT 170.6950 64.6650 172.6950 66.6650 ;
        RECT 162.1800 64.6650 164.1800 66.6650 ;
        RECT 153.6650 64.6650 155.6650 66.6650 ;
        RECT 145.1500 64.6650 147.1500 66.6650 ;
        RECT 255.8450 64.6650 257.8450 66.6650 ;
        RECT 247.3300 64.6650 249.3300 66.6650 ;
        RECT 238.8150 64.6650 240.8150 66.6650 ;
        RECT 230.3000 64.6650 232.3000 66.6650 ;
        RECT 221.7850 64.6650 223.7850 66.6650 ;
        RECT 213.2700 64.6650 215.2700 66.6650 ;
        RECT 264.3600 64.6650 266.3600 66.6650 ;
        RECT 272.8750 64.6650 274.8750 66.6650 ;
        RECT 145.1500 85.9500 147.1500 87.9500 ;
        RECT 153.6650 85.9500 155.6650 87.9500 ;
        RECT 162.1800 85.9500 164.1800 87.9500 ;
        RECT 170.6950 85.9500 172.6950 87.9500 ;
        RECT 170.6950 78.8550 172.6950 80.8550 ;
        RECT 162.1800 78.8550 164.1800 80.8550 ;
        RECT 153.6650 78.8550 155.6650 80.8550 ;
        RECT 145.1500 78.8550 147.1500 80.8550 ;
        RECT 170.6950 71.7600 172.6950 73.7600 ;
        RECT 162.1800 71.7600 164.1800 73.7600 ;
        RECT 153.6650 71.7600 155.6650 73.7600 ;
        RECT 145.1500 71.7600 147.1500 73.7600 ;
        RECT 145.1500 93.0450 147.1500 95.0450 ;
        RECT 153.6650 93.0450 155.6650 95.0450 ;
        RECT 162.1800 93.0450 164.1800 95.0450 ;
        RECT 170.6950 93.0450 172.6950 95.0450 ;
        RECT 145.1500 100.1400 147.1500 102.1400 ;
        RECT 153.6650 100.1400 155.6650 102.1400 ;
        RECT 162.1800 100.1400 164.1800 102.1400 ;
        RECT 170.6950 100.1400 172.6950 102.1400 ;
        RECT 179.2100 85.9500 181.2100 87.9500 ;
        RECT 187.7250 85.9500 189.7250 87.9500 ;
        RECT 196.2400 85.9500 198.2400 87.9500 ;
        RECT 204.7550 85.9500 206.7550 87.9500 ;
        RECT 204.7550 78.8550 206.7550 80.8550 ;
        RECT 196.2400 78.8550 198.2400 80.8550 ;
        RECT 187.7250 78.8550 189.7250 80.8550 ;
        RECT 179.2100 78.8550 181.2100 80.8550 ;
        RECT 204.7550 71.7600 206.7550 73.7600 ;
        RECT 196.2400 71.7600 198.2400 73.7600 ;
        RECT 187.7250 71.7600 189.7250 73.7600 ;
        RECT 179.2100 71.7600 181.2100 73.7600 ;
        RECT 179.2100 93.0450 181.2100 95.0450 ;
        RECT 187.7250 93.0450 189.7250 95.0450 ;
        RECT 196.2400 93.0450 198.2400 95.0450 ;
        RECT 204.7550 93.0450 206.7550 95.0450 ;
        RECT 179.2100 100.1400 181.2100 102.1400 ;
        RECT 187.7250 100.1400 189.7250 102.1400 ;
        RECT 196.2400 100.1400 198.2400 102.1400 ;
        RECT 204.7550 100.1400 206.7550 102.1400 ;
        RECT 145.1500 121.4250 147.1500 123.4250 ;
        RECT 153.6650 121.4250 155.6650 123.4250 ;
        RECT 162.1800 121.4250 164.1800 123.4250 ;
        RECT 170.6950 121.4250 172.6950 123.4250 ;
        RECT 170.6950 114.3300 172.6950 116.3300 ;
        RECT 162.1800 114.3300 164.1800 116.3300 ;
        RECT 153.6650 114.3300 155.6650 116.3300 ;
        RECT 145.1500 114.3300 147.1500 116.3300 ;
        RECT 170.6950 107.2350 172.6950 109.2350 ;
        RECT 162.1800 107.2350 164.1800 109.2350 ;
        RECT 153.6650 107.2350 155.6650 109.2350 ;
        RECT 145.1500 107.2350 147.1500 109.2350 ;
        RECT 145.1500 128.5200 147.1500 130.5200 ;
        RECT 153.6650 128.5200 155.6650 130.5200 ;
        RECT 162.1800 128.5200 164.1800 130.5200 ;
        RECT 170.6950 128.5200 172.6950 130.5200 ;
        RECT 145.1500 135.6150 147.1500 137.6150 ;
        RECT 153.6650 135.6150 155.6650 137.6150 ;
        RECT 162.1800 135.6150 164.1800 137.6150 ;
        RECT 170.6950 135.6150 172.6950 137.6150 ;
        RECT 179.2100 121.4250 181.2100 123.4250 ;
        RECT 187.7250 121.4250 189.7250 123.4250 ;
        RECT 196.2400 121.4250 198.2400 123.4250 ;
        RECT 204.7550 121.4250 206.7550 123.4250 ;
        RECT 204.7550 114.3300 206.7550 116.3300 ;
        RECT 196.2400 114.3300 198.2400 116.3300 ;
        RECT 187.7250 114.3300 189.7250 116.3300 ;
        RECT 179.2100 114.3300 181.2100 116.3300 ;
        RECT 204.7550 107.2350 206.7550 109.2350 ;
        RECT 196.2400 107.2350 198.2400 109.2350 ;
        RECT 187.7250 107.2350 189.7250 109.2350 ;
        RECT 179.2100 107.2350 181.2100 109.2350 ;
        RECT 179.2100 128.5200 181.2100 130.5200 ;
        RECT 187.7250 128.5200 189.7250 130.5200 ;
        RECT 196.2400 128.5200 198.2400 130.5200 ;
        RECT 204.7550 128.5200 206.7550 130.5200 ;
        RECT 179.2100 135.6150 181.2100 137.6150 ;
        RECT 187.7250 135.6150 189.7250 137.6150 ;
        RECT 196.2400 135.6150 198.2400 137.6150 ;
        RECT 204.7550 135.6150 206.7550 137.6150 ;
        RECT 213.2700 85.9500 215.2700 87.9500 ;
        RECT 221.7850 85.9500 223.7850 87.9500 ;
        RECT 230.3000 85.9500 232.3000 87.9500 ;
        RECT 238.8150 85.9500 240.8150 87.9500 ;
        RECT 238.8150 78.8550 240.8150 80.8550 ;
        RECT 230.3000 78.8550 232.3000 80.8550 ;
        RECT 221.7850 78.8550 223.7850 80.8550 ;
        RECT 213.2700 78.8550 215.2700 80.8550 ;
        RECT 238.8150 71.7600 240.8150 73.7600 ;
        RECT 230.3000 71.7600 232.3000 73.7600 ;
        RECT 221.7850 71.7600 223.7850 73.7600 ;
        RECT 213.2700 71.7600 215.2700 73.7600 ;
        RECT 213.2700 93.0450 215.2700 95.0450 ;
        RECT 221.7850 93.0450 223.7850 95.0450 ;
        RECT 230.3000 93.0450 232.3000 95.0450 ;
        RECT 238.8150 93.0450 240.8150 95.0450 ;
        RECT 213.2700 100.1400 215.2700 102.1400 ;
        RECT 221.7850 100.1400 223.7850 102.1400 ;
        RECT 230.3000 100.1400 232.3000 102.1400 ;
        RECT 238.8150 100.1400 240.8150 102.1400 ;
        RECT 247.3300 85.9500 249.3300 87.9500 ;
        RECT 255.8450 85.9500 257.8450 87.9500 ;
        RECT 264.3600 85.9500 266.3600 87.9500 ;
        RECT 272.8750 85.9500 274.8750 87.9500 ;
        RECT 272.8750 78.8550 274.8750 80.8550 ;
        RECT 264.3600 78.8550 266.3600 80.8550 ;
        RECT 255.8450 78.8550 257.8450 80.8550 ;
        RECT 247.3300 78.8550 249.3300 80.8550 ;
        RECT 272.8750 71.7600 274.8750 73.7600 ;
        RECT 264.3600 71.7600 266.3600 73.7600 ;
        RECT 255.8450 71.7600 257.8450 73.7600 ;
        RECT 247.3300 71.7600 249.3300 73.7600 ;
        RECT 247.3300 93.0450 249.3300 95.0450 ;
        RECT 255.8450 93.0450 257.8450 95.0450 ;
        RECT 264.3600 93.0450 266.3600 95.0450 ;
        RECT 272.8750 93.0450 274.8750 95.0450 ;
        RECT 247.3300 100.1400 249.3300 102.1400 ;
        RECT 255.8450 100.1400 257.8450 102.1400 ;
        RECT 264.3600 100.1400 266.3600 102.1400 ;
        RECT 272.8750 100.1400 274.8750 102.1400 ;
        RECT 213.2700 121.4250 215.2700 123.4250 ;
        RECT 221.7850 121.4250 223.7850 123.4250 ;
        RECT 230.3000 121.4250 232.3000 123.4250 ;
        RECT 238.8150 121.4250 240.8150 123.4250 ;
        RECT 238.8150 114.3300 240.8150 116.3300 ;
        RECT 230.3000 114.3300 232.3000 116.3300 ;
        RECT 221.7850 114.3300 223.7850 116.3300 ;
        RECT 213.2700 114.3300 215.2700 116.3300 ;
        RECT 238.8150 107.2350 240.8150 109.2350 ;
        RECT 230.3000 107.2350 232.3000 109.2350 ;
        RECT 221.7850 107.2350 223.7850 109.2350 ;
        RECT 213.2700 107.2350 215.2700 109.2350 ;
        RECT 213.2700 128.5200 215.2700 130.5200 ;
        RECT 221.7850 128.5200 223.7850 130.5200 ;
        RECT 230.3000 128.5200 232.3000 130.5200 ;
        RECT 238.8150 128.5200 240.8150 130.5200 ;
        RECT 213.2700 135.6150 215.2700 137.6150 ;
        RECT 221.7850 135.6150 223.7850 137.6150 ;
        RECT 230.3000 135.6150 232.3000 137.6150 ;
        RECT 238.8150 135.6150 240.8150 137.6150 ;
        RECT 247.3300 121.4250 249.3300 123.4250 ;
        RECT 255.8450 121.4250 257.8450 123.4250 ;
        RECT 264.3600 121.4250 266.3600 123.4250 ;
        RECT 272.8750 121.4250 274.8750 123.4250 ;
        RECT 272.8750 114.3300 274.8750 116.3300 ;
        RECT 264.3600 114.3300 266.3600 116.3300 ;
        RECT 255.8450 114.3300 257.8450 116.3300 ;
        RECT 247.3300 114.3300 249.3300 116.3300 ;
        RECT 272.8750 107.2350 274.8750 109.2350 ;
        RECT 264.3600 107.2350 266.3600 109.2350 ;
        RECT 255.8450 107.2350 257.8450 109.2350 ;
        RECT 247.3300 107.2350 249.3300 109.2350 ;
        RECT 247.3300 128.5200 249.3300 130.5200 ;
        RECT 255.8450 128.5200 257.8450 130.5200 ;
        RECT 264.3600 128.5200 266.3600 130.5200 ;
        RECT 272.8750 128.5200 274.8750 130.5200 ;
        RECT 247.3300 135.6150 249.3300 137.6150 ;
        RECT 255.8450 135.6150 257.8450 137.6150 ;
        RECT 264.3600 135.6150 266.3600 137.6150 ;
        RECT 272.8750 135.6150 274.8750 137.6150 ;
        RECT 68.5150 142.7100 70.5150 144.7100 ;
        RECT 68.5150 149.8050 70.5150 151.8050 ;
        RECT 68.5150 156.9000 70.5150 158.9000 ;
        RECT 68.5150 163.9950 70.5150 165.9950 ;
        RECT 68.5150 171.0900 70.5150 173.0900 ;
        RECT 68.5150 178.1850 70.5150 180.1850 ;
        RECT 68.5150 185.2800 70.5150 187.2800 ;
        RECT 68.5150 192.3750 70.5150 194.3750 ;
        RECT 68.5150 199.4700 70.5150 201.4700 ;
        RECT 68.5150 206.5650 70.5150 208.5650 ;
        RECT 6.0000 156.9000 8.0000 158.9000 ;
        RECT 6.0000 149.8050 8.0000 151.8050 ;
        RECT 6.0000 142.7100 8.0000 144.7100 ;
        RECT 6.0000 171.0900 8.0000 173.0900 ;
        RECT 6.0000 163.9950 8.0000 165.9950 ;
        RECT 44.0000 156.9000 46.0000 158.9000 ;
        RECT 60.0000 156.9000 62.0000 158.9000 ;
        RECT 44.0000 149.8050 46.0000 151.8050 ;
        RECT 44.0000 142.7100 46.0000 144.7100 ;
        RECT 60.0000 142.7100 62.0000 144.7100 ;
        RECT 60.0000 149.8050 62.0000 151.8050 ;
        RECT 44.0000 171.0900 46.0000 173.0900 ;
        RECT 44.0000 163.9950 46.0000 165.9950 ;
        RECT 60.0000 163.9950 62.0000 165.9950 ;
        RECT 60.0000 171.0900 62.0000 173.0900 ;
        RECT 6.0000 192.3750 8.0000 194.3750 ;
        RECT 6.0000 178.1850 8.0000 180.1850 ;
        RECT 6.0000 185.2800 8.0000 187.2800 ;
        RECT 6.0000 199.4700 8.0000 201.4700 ;
        RECT 6.0000 206.5650 8.0000 208.5650 ;
        RECT 44.0000 192.3750 46.0000 194.3750 ;
        RECT 60.0000 192.3750 62.0000 194.3750 ;
        RECT 44.0000 178.1850 46.0000 180.1850 ;
        RECT 44.0000 185.2800 46.0000 187.2800 ;
        RECT 60.0000 185.2800 62.0000 187.2800 ;
        RECT 60.0000 178.1850 62.0000 180.1850 ;
        RECT 44.0000 199.4700 46.0000 201.4700 ;
        RECT 44.0000 206.5650 46.0000 208.5650 ;
        RECT 60.0000 206.5650 62.0000 208.5650 ;
        RECT 60.0000 199.4700 62.0000 201.4700 ;
        RECT 77.0300 156.9000 79.0300 158.9000 ;
        RECT 85.5450 156.9000 87.5450 158.9000 ;
        RECT 94.0600 156.9000 96.0600 158.9000 ;
        RECT 102.5750 156.9000 104.5750 158.9000 ;
        RECT 102.5750 149.8050 104.5750 151.8050 ;
        RECT 94.0600 149.8050 96.0600 151.8050 ;
        RECT 85.5450 149.8050 87.5450 151.8050 ;
        RECT 77.0300 149.8050 79.0300 151.8050 ;
        RECT 102.5750 142.7100 104.5750 144.7100 ;
        RECT 94.0600 142.7100 96.0600 144.7100 ;
        RECT 85.5450 142.7100 87.5450 144.7100 ;
        RECT 77.0300 142.7100 79.0300 144.7100 ;
        RECT 77.0300 163.9950 79.0300 165.9950 ;
        RECT 85.5450 163.9950 87.5450 165.9950 ;
        RECT 94.0600 163.9950 96.0600 165.9950 ;
        RECT 102.5750 163.9950 104.5750 165.9950 ;
        RECT 77.0300 171.0900 79.0300 173.0900 ;
        RECT 85.5450 171.0900 87.5450 173.0900 ;
        RECT 94.0600 171.0900 96.0600 173.0900 ;
        RECT 102.5750 171.0900 104.5750 173.0900 ;
        RECT 111.0900 156.9000 113.0900 158.9000 ;
        RECT 119.6050 156.9000 121.6050 158.9000 ;
        RECT 128.1200 156.9000 130.1200 158.9000 ;
        RECT 136.6350 156.9000 138.6350 158.9000 ;
        RECT 136.6350 149.8050 138.6350 151.8050 ;
        RECT 128.1200 149.8050 130.1200 151.8050 ;
        RECT 119.6050 149.8050 121.6050 151.8050 ;
        RECT 111.0900 149.8050 113.0900 151.8050 ;
        RECT 136.6350 142.7100 138.6350 144.7100 ;
        RECT 128.1200 142.7100 130.1200 144.7100 ;
        RECT 119.6050 142.7100 121.6050 144.7100 ;
        RECT 111.0900 142.7100 113.0900 144.7100 ;
        RECT 111.0900 163.9950 113.0900 165.9950 ;
        RECT 119.6050 163.9950 121.6050 165.9950 ;
        RECT 128.1200 163.9950 130.1200 165.9950 ;
        RECT 136.6350 163.9950 138.6350 165.9950 ;
        RECT 111.0900 171.0900 113.0900 173.0900 ;
        RECT 119.6050 171.0900 121.6050 173.0900 ;
        RECT 128.1200 171.0900 130.1200 173.0900 ;
        RECT 136.6350 171.0900 138.6350 173.0900 ;
        RECT 77.0300 192.3750 79.0300 194.3750 ;
        RECT 85.5450 192.3750 87.5450 194.3750 ;
        RECT 94.0600 192.3750 96.0600 194.3750 ;
        RECT 102.5750 192.3750 104.5750 194.3750 ;
        RECT 102.5750 185.2800 104.5750 187.2800 ;
        RECT 94.0600 185.2800 96.0600 187.2800 ;
        RECT 85.5450 185.2800 87.5450 187.2800 ;
        RECT 77.0300 185.2800 79.0300 187.2800 ;
        RECT 102.5750 178.1850 104.5750 180.1850 ;
        RECT 94.0600 178.1850 96.0600 180.1850 ;
        RECT 85.5450 178.1850 87.5450 180.1850 ;
        RECT 77.0300 178.1850 79.0300 180.1850 ;
        RECT 77.0300 199.4700 79.0300 201.4700 ;
        RECT 85.5450 199.4700 87.5450 201.4700 ;
        RECT 94.0600 199.4700 96.0600 201.4700 ;
        RECT 102.5750 199.4700 104.5750 201.4700 ;
        RECT 77.0300 206.5650 79.0300 208.5650 ;
        RECT 85.5450 206.5650 87.5450 208.5650 ;
        RECT 94.0600 206.5650 96.0600 208.5650 ;
        RECT 102.5750 206.5650 104.5750 208.5650 ;
        RECT 111.0900 192.3750 113.0900 194.3750 ;
        RECT 119.6050 192.3750 121.6050 194.3750 ;
        RECT 128.1200 192.3750 130.1200 194.3750 ;
        RECT 136.6350 192.3750 138.6350 194.3750 ;
        RECT 136.6350 185.2800 138.6350 187.2800 ;
        RECT 128.1200 185.2800 130.1200 187.2800 ;
        RECT 119.6050 185.2800 121.6050 187.2800 ;
        RECT 111.0900 185.2800 113.0900 187.2800 ;
        RECT 136.6350 178.1850 138.6350 180.1850 ;
        RECT 128.1200 178.1850 130.1200 180.1850 ;
        RECT 119.6050 178.1850 121.6050 180.1850 ;
        RECT 111.0900 178.1850 113.0900 180.1850 ;
        RECT 111.0900 199.4700 113.0900 201.4700 ;
        RECT 119.6050 199.4700 121.6050 201.4700 ;
        RECT 128.1200 199.4700 130.1200 201.4700 ;
        RECT 136.6350 199.4700 138.6350 201.4700 ;
        RECT 111.0900 206.5650 113.0900 208.5650 ;
        RECT 119.6050 206.5650 121.6050 208.5650 ;
        RECT 128.1200 206.5650 130.1200 208.5650 ;
        RECT 136.6350 206.5650 138.6350 208.5650 ;
        RECT 68.5150 213.6600 70.5150 215.6600 ;
        RECT 68.5150 220.7550 70.5150 222.7550 ;
        RECT 68.5150 227.8500 70.5150 229.8500 ;
        RECT 68.5150 234.9450 70.5150 236.9450 ;
        RECT 68.5150 242.0400 70.5150 244.0400 ;
        RECT 68.5150 249.1350 70.5150 251.1350 ;
        RECT 68.5150 256.2300 70.5150 258.2300 ;
        RECT 68.5150 263.3250 70.5150 265.3250 ;
        RECT 68.5150 270.4200 70.5150 272.4200 ;
        RECT 68.5150 277.5150 70.5150 279.5150 ;
        RECT 6.0000 220.7550 8.0000 222.7550 ;
        RECT 6.0000 213.6600 8.0000 215.6600 ;
        RECT 6.0000 234.9450 8.0000 236.9450 ;
        RECT 6.0000 227.8500 8.0000 229.8500 ;
        RECT 6.0000 242.0400 8.0000 244.0400 ;
        RECT 44.0000 220.7550 46.0000 222.7550 ;
        RECT 44.0000 213.6600 46.0000 215.6600 ;
        RECT 60.0000 213.6600 62.0000 215.6600 ;
        RECT 60.0000 220.7550 62.0000 222.7550 ;
        RECT 44.0000 227.8500 46.0000 229.8500 ;
        RECT 44.0000 234.9450 46.0000 236.9450 ;
        RECT 44.0000 242.0400 46.0000 244.0400 ;
        RECT 60.0000 227.8500 62.0000 229.8500 ;
        RECT 60.0000 234.9450 62.0000 236.9450 ;
        RECT 60.0000 242.0400 62.0000 244.0400 ;
        RECT 6.0000 249.1350 8.0000 251.1350 ;
        RECT 6.0000 256.2300 8.0000 258.2300 ;
        RECT 6.0000 270.4200 8.0000 272.4200 ;
        RECT 6.0000 263.3250 8.0000 265.3250 ;
        RECT 6.0000 277.5150 8.0000 279.5150 ;
        RECT 44.0000 249.1350 46.0000 251.1350 ;
        RECT 44.0000 256.2300 46.0000 258.2300 ;
        RECT 60.0000 256.2300 62.0000 258.2300 ;
        RECT 60.0000 249.1350 62.0000 251.1350 ;
        RECT 44.0000 263.3250 46.0000 265.3250 ;
        RECT 44.0000 270.4200 46.0000 272.4200 ;
        RECT 44.0000 277.5150 46.0000 279.5150 ;
        RECT 60.0000 270.4200 62.0000 272.4200 ;
        RECT 60.0000 263.3250 62.0000 265.3250 ;
        RECT 60.0000 277.5150 62.0000 279.5150 ;
        RECT 102.5750 220.7550 104.5750 222.7550 ;
        RECT 94.0600 220.7550 96.0600 222.7550 ;
        RECT 85.5450 220.7550 87.5450 222.7550 ;
        RECT 77.0300 220.7550 79.0300 222.7550 ;
        RECT 102.5750 213.6600 104.5750 215.6600 ;
        RECT 94.0600 213.6600 96.0600 215.6600 ;
        RECT 85.5450 213.6600 87.5450 215.6600 ;
        RECT 77.0300 213.6600 79.0300 215.6600 ;
        RECT 85.5450 227.8500 87.5450 229.8500 ;
        RECT 77.0300 227.8500 79.0300 229.8500 ;
        RECT 94.0600 227.8500 96.0600 229.8500 ;
        RECT 102.5750 227.8500 104.5750 229.8500 ;
        RECT 77.0300 234.9450 79.0300 236.9450 ;
        RECT 85.5450 234.9450 87.5450 236.9450 ;
        RECT 94.0600 234.9450 96.0600 236.9450 ;
        RECT 102.5750 234.9450 104.5750 236.9450 ;
        RECT 77.0300 242.0400 79.0300 244.0400 ;
        RECT 85.5450 242.0400 87.5450 244.0400 ;
        RECT 94.0600 242.0400 96.0600 244.0400 ;
        RECT 102.5750 242.0400 104.5750 244.0400 ;
        RECT 136.6350 220.7550 138.6350 222.7550 ;
        RECT 128.1200 220.7550 130.1200 222.7550 ;
        RECT 119.6050 220.7550 121.6050 222.7550 ;
        RECT 111.0900 220.7550 113.0900 222.7550 ;
        RECT 136.6350 213.6600 138.6350 215.6600 ;
        RECT 128.1200 213.6600 130.1200 215.6600 ;
        RECT 119.6050 213.6600 121.6050 215.6600 ;
        RECT 111.0900 213.6600 113.0900 215.6600 ;
        RECT 119.6050 227.8500 121.6050 229.8500 ;
        RECT 111.0900 227.8500 113.0900 229.8500 ;
        RECT 128.1200 227.8500 130.1200 229.8500 ;
        RECT 136.6350 227.8500 138.6350 229.8500 ;
        RECT 111.0900 234.9450 113.0900 236.9450 ;
        RECT 119.6050 234.9450 121.6050 236.9450 ;
        RECT 128.1200 234.9450 130.1200 236.9450 ;
        RECT 136.6350 234.9450 138.6350 236.9450 ;
        RECT 111.0900 242.0400 113.0900 244.0400 ;
        RECT 119.6050 242.0400 121.6050 244.0400 ;
        RECT 128.1200 242.0400 130.1200 244.0400 ;
        RECT 136.6350 242.0400 138.6350 244.0400 ;
        RECT 102.5750 256.2300 104.5750 258.2300 ;
        RECT 94.0600 256.2300 96.0600 258.2300 ;
        RECT 85.5450 256.2300 87.5450 258.2300 ;
        RECT 77.0300 256.2300 79.0300 258.2300 ;
        RECT 102.5750 249.1350 104.5750 251.1350 ;
        RECT 94.0600 249.1350 96.0600 251.1350 ;
        RECT 85.5450 249.1350 87.5450 251.1350 ;
        RECT 77.0300 249.1350 79.0300 251.1350 ;
        RECT 85.5450 263.3250 87.5450 265.3250 ;
        RECT 77.0300 263.3250 79.0300 265.3250 ;
        RECT 94.0600 263.3250 96.0600 265.3250 ;
        RECT 102.5750 263.3250 104.5750 265.3250 ;
        RECT 77.0300 270.4200 79.0300 272.4200 ;
        RECT 85.5450 270.4200 87.5450 272.4200 ;
        RECT 94.0600 270.4200 96.0600 272.4200 ;
        RECT 102.5750 270.4200 104.5750 272.4200 ;
        RECT 77.0300 277.5150 79.0300 279.5150 ;
        RECT 85.5450 277.5150 87.5450 279.5150 ;
        RECT 94.0600 277.5150 96.0600 279.5150 ;
        RECT 102.5750 277.5150 104.5750 279.5150 ;
        RECT 136.6350 256.2300 138.6350 258.2300 ;
        RECT 128.1200 256.2300 130.1200 258.2300 ;
        RECT 119.6050 256.2300 121.6050 258.2300 ;
        RECT 111.0900 256.2300 113.0900 258.2300 ;
        RECT 136.6350 249.1350 138.6350 251.1350 ;
        RECT 128.1200 249.1350 130.1200 251.1350 ;
        RECT 119.6050 249.1350 121.6050 251.1350 ;
        RECT 111.0900 249.1350 113.0900 251.1350 ;
        RECT 119.6050 263.3250 121.6050 265.3250 ;
        RECT 111.0900 263.3250 113.0900 265.3250 ;
        RECT 128.1200 263.3250 130.1200 265.3250 ;
        RECT 136.6350 263.3250 138.6350 265.3250 ;
        RECT 111.0900 270.4200 113.0900 272.4200 ;
        RECT 119.6050 270.4200 121.6050 272.4200 ;
        RECT 128.1200 270.4200 130.1200 272.4200 ;
        RECT 136.6350 270.4200 138.6350 272.4200 ;
        RECT 111.0900 277.5150 113.0900 279.5150 ;
        RECT 119.6050 277.5150 121.6050 279.5150 ;
        RECT 128.1200 277.5150 130.1200 279.5150 ;
        RECT 136.6350 277.5150 138.6350 279.5150 ;
        RECT 145.1500 156.9000 147.1500 158.9000 ;
        RECT 153.6650 156.9000 155.6650 158.9000 ;
        RECT 162.1800 156.9000 164.1800 158.9000 ;
        RECT 170.6950 156.9000 172.6950 158.9000 ;
        RECT 170.6950 149.8050 172.6950 151.8050 ;
        RECT 162.1800 149.8050 164.1800 151.8050 ;
        RECT 153.6650 149.8050 155.6650 151.8050 ;
        RECT 145.1500 149.8050 147.1500 151.8050 ;
        RECT 170.6950 142.7100 172.6950 144.7100 ;
        RECT 162.1800 142.7100 164.1800 144.7100 ;
        RECT 153.6650 142.7100 155.6650 144.7100 ;
        RECT 145.1500 142.7100 147.1500 144.7100 ;
        RECT 145.1500 163.9950 147.1500 165.9950 ;
        RECT 153.6650 163.9950 155.6650 165.9950 ;
        RECT 162.1800 163.9950 164.1800 165.9950 ;
        RECT 170.6950 163.9950 172.6950 165.9950 ;
        RECT 145.1500 171.0900 147.1500 173.0900 ;
        RECT 153.6650 171.0900 155.6650 173.0900 ;
        RECT 162.1800 171.0900 164.1800 173.0900 ;
        RECT 170.6950 171.0900 172.6950 173.0900 ;
        RECT 179.2100 156.9000 181.2100 158.9000 ;
        RECT 187.7250 156.9000 189.7250 158.9000 ;
        RECT 196.2400 156.9000 198.2400 158.9000 ;
        RECT 204.7550 156.9000 206.7550 158.9000 ;
        RECT 204.7550 149.8050 206.7550 151.8050 ;
        RECT 196.2400 149.8050 198.2400 151.8050 ;
        RECT 187.7250 149.8050 189.7250 151.8050 ;
        RECT 179.2100 149.8050 181.2100 151.8050 ;
        RECT 204.7550 142.7100 206.7550 144.7100 ;
        RECT 196.2400 142.7100 198.2400 144.7100 ;
        RECT 187.7250 142.7100 189.7250 144.7100 ;
        RECT 179.2100 142.7100 181.2100 144.7100 ;
        RECT 179.2100 163.9950 181.2100 165.9950 ;
        RECT 187.7250 163.9950 189.7250 165.9950 ;
        RECT 196.2400 163.9950 198.2400 165.9950 ;
        RECT 204.7550 163.9950 206.7550 165.9950 ;
        RECT 179.2100 171.0900 181.2100 173.0900 ;
        RECT 187.7250 171.0900 189.7250 173.0900 ;
        RECT 196.2400 171.0900 198.2400 173.0900 ;
        RECT 204.7550 171.0900 206.7550 173.0900 ;
        RECT 145.1500 192.3750 147.1500 194.3750 ;
        RECT 153.6650 192.3750 155.6650 194.3750 ;
        RECT 162.1800 192.3750 164.1800 194.3750 ;
        RECT 170.6950 192.3750 172.6950 194.3750 ;
        RECT 170.6950 185.2800 172.6950 187.2800 ;
        RECT 162.1800 185.2800 164.1800 187.2800 ;
        RECT 153.6650 185.2800 155.6650 187.2800 ;
        RECT 145.1500 185.2800 147.1500 187.2800 ;
        RECT 170.6950 178.1850 172.6950 180.1850 ;
        RECT 162.1800 178.1850 164.1800 180.1850 ;
        RECT 153.6650 178.1850 155.6650 180.1850 ;
        RECT 145.1500 178.1850 147.1500 180.1850 ;
        RECT 145.1500 199.4700 147.1500 201.4700 ;
        RECT 153.6650 199.4700 155.6650 201.4700 ;
        RECT 162.1800 199.4700 164.1800 201.4700 ;
        RECT 170.6950 199.4700 172.6950 201.4700 ;
        RECT 145.1500 206.5650 147.1500 208.5650 ;
        RECT 153.6650 206.5650 155.6650 208.5650 ;
        RECT 162.1800 206.5650 164.1800 208.5650 ;
        RECT 170.6950 206.5650 172.6950 208.5650 ;
        RECT 179.2100 192.3750 181.2100 194.3750 ;
        RECT 187.7250 192.3750 189.7250 194.3750 ;
        RECT 196.2400 192.3750 198.2400 194.3750 ;
        RECT 204.7550 192.3750 206.7550 194.3750 ;
        RECT 204.7550 185.2800 206.7550 187.2800 ;
        RECT 196.2400 185.2800 198.2400 187.2800 ;
        RECT 187.7250 185.2800 189.7250 187.2800 ;
        RECT 179.2100 185.2800 181.2100 187.2800 ;
        RECT 204.7550 178.1850 206.7550 180.1850 ;
        RECT 196.2400 178.1850 198.2400 180.1850 ;
        RECT 187.7250 178.1850 189.7250 180.1850 ;
        RECT 179.2100 178.1850 181.2100 180.1850 ;
        RECT 179.2100 199.4700 181.2100 201.4700 ;
        RECT 187.7250 199.4700 189.7250 201.4700 ;
        RECT 196.2400 199.4700 198.2400 201.4700 ;
        RECT 204.7550 199.4700 206.7550 201.4700 ;
        RECT 179.2100 206.5650 181.2100 208.5650 ;
        RECT 187.7250 206.5650 189.7250 208.5650 ;
        RECT 196.2400 206.5650 198.2400 208.5650 ;
        RECT 204.7550 206.5650 206.7550 208.5650 ;
        RECT 213.2700 156.9000 215.2700 158.9000 ;
        RECT 221.7850 156.9000 223.7850 158.9000 ;
        RECT 230.3000 156.9000 232.3000 158.9000 ;
        RECT 238.8150 156.9000 240.8150 158.9000 ;
        RECT 238.8150 149.8050 240.8150 151.8050 ;
        RECT 230.3000 149.8050 232.3000 151.8050 ;
        RECT 221.7850 149.8050 223.7850 151.8050 ;
        RECT 213.2700 149.8050 215.2700 151.8050 ;
        RECT 238.8150 142.7100 240.8150 144.7100 ;
        RECT 230.3000 142.7100 232.3000 144.7100 ;
        RECT 221.7850 142.7100 223.7850 144.7100 ;
        RECT 213.2700 142.7100 215.2700 144.7100 ;
        RECT 213.2700 163.9950 215.2700 165.9950 ;
        RECT 221.7850 163.9950 223.7850 165.9950 ;
        RECT 230.3000 163.9950 232.3000 165.9950 ;
        RECT 238.8150 163.9950 240.8150 165.9950 ;
        RECT 213.2700 171.0900 215.2700 173.0900 ;
        RECT 221.7850 171.0900 223.7850 173.0900 ;
        RECT 230.3000 171.0900 232.3000 173.0900 ;
        RECT 238.8150 171.0900 240.8150 173.0900 ;
        RECT 247.3300 156.9000 249.3300 158.9000 ;
        RECT 255.8450 156.9000 257.8450 158.9000 ;
        RECT 264.3600 156.9000 266.3600 158.9000 ;
        RECT 272.8750 156.9000 274.8750 158.9000 ;
        RECT 272.8750 149.8050 274.8750 151.8050 ;
        RECT 264.3600 149.8050 266.3600 151.8050 ;
        RECT 255.8450 149.8050 257.8450 151.8050 ;
        RECT 247.3300 149.8050 249.3300 151.8050 ;
        RECT 272.8750 142.7100 274.8750 144.7100 ;
        RECT 264.3600 142.7100 266.3600 144.7100 ;
        RECT 255.8450 142.7100 257.8450 144.7100 ;
        RECT 247.3300 142.7100 249.3300 144.7100 ;
        RECT 247.3300 163.9950 249.3300 165.9950 ;
        RECT 255.8450 163.9950 257.8450 165.9950 ;
        RECT 264.3600 163.9950 266.3600 165.9950 ;
        RECT 272.8750 163.9950 274.8750 165.9950 ;
        RECT 247.3300 171.0900 249.3300 173.0900 ;
        RECT 255.8450 171.0900 257.8450 173.0900 ;
        RECT 264.3600 171.0900 266.3600 173.0900 ;
        RECT 272.8750 171.0900 274.8750 173.0900 ;
        RECT 213.2700 192.3750 215.2700 194.3750 ;
        RECT 221.7850 192.3750 223.7850 194.3750 ;
        RECT 230.3000 192.3750 232.3000 194.3750 ;
        RECT 238.8150 192.3750 240.8150 194.3750 ;
        RECT 238.8150 185.2800 240.8150 187.2800 ;
        RECT 230.3000 185.2800 232.3000 187.2800 ;
        RECT 221.7850 185.2800 223.7850 187.2800 ;
        RECT 213.2700 185.2800 215.2700 187.2800 ;
        RECT 238.8150 178.1850 240.8150 180.1850 ;
        RECT 230.3000 178.1850 232.3000 180.1850 ;
        RECT 221.7850 178.1850 223.7850 180.1850 ;
        RECT 213.2700 178.1850 215.2700 180.1850 ;
        RECT 213.2700 199.4700 215.2700 201.4700 ;
        RECT 221.7850 199.4700 223.7850 201.4700 ;
        RECT 230.3000 199.4700 232.3000 201.4700 ;
        RECT 238.8150 199.4700 240.8150 201.4700 ;
        RECT 213.2700 206.5650 215.2700 208.5650 ;
        RECT 221.7850 206.5650 223.7850 208.5650 ;
        RECT 230.3000 206.5650 232.3000 208.5650 ;
        RECT 238.8150 206.5650 240.8150 208.5650 ;
        RECT 247.3300 192.3750 249.3300 194.3750 ;
        RECT 255.8450 192.3750 257.8450 194.3750 ;
        RECT 264.3600 192.3750 266.3600 194.3750 ;
        RECT 272.8750 192.3750 274.8750 194.3750 ;
        RECT 272.8750 185.2800 274.8750 187.2800 ;
        RECT 264.3600 185.2800 266.3600 187.2800 ;
        RECT 255.8450 185.2800 257.8450 187.2800 ;
        RECT 247.3300 185.2800 249.3300 187.2800 ;
        RECT 272.8750 178.1850 274.8750 180.1850 ;
        RECT 264.3600 178.1850 266.3600 180.1850 ;
        RECT 255.8450 178.1850 257.8450 180.1850 ;
        RECT 247.3300 178.1850 249.3300 180.1850 ;
        RECT 247.3300 199.4700 249.3300 201.4700 ;
        RECT 255.8450 199.4700 257.8450 201.4700 ;
        RECT 264.3600 199.4700 266.3600 201.4700 ;
        RECT 272.8750 199.4700 274.8750 201.4700 ;
        RECT 247.3300 206.5650 249.3300 208.5650 ;
        RECT 255.8450 206.5650 257.8450 208.5650 ;
        RECT 264.3600 206.5650 266.3600 208.5650 ;
        RECT 272.8750 206.5650 274.8750 208.5650 ;
        RECT 170.6950 220.7550 172.6950 222.7550 ;
        RECT 162.1800 220.7550 164.1800 222.7550 ;
        RECT 153.6650 220.7550 155.6650 222.7550 ;
        RECT 145.1500 220.7550 147.1500 222.7550 ;
        RECT 170.6950 213.6600 172.6950 215.6600 ;
        RECT 162.1800 213.6600 164.1800 215.6600 ;
        RECT 153.6650 213.6600 155.6650 215.6600 ;
        RECT 145.1500 213.6600 147.1500 215.6600 ;
        RECT 153.6650 227.8500 155.6650 229.8500 ;
        RECT 145.1500 227.8500 147.1500 229.8500 ;
        RECT 162.1800 227.8500 164.1800 229.8500 ;
        RECT 170.6950 227.8500 172.6950 229.8500 ;
        RECT 145.1500 234.9450 147.1500 236.9450 ;
        RECT 153.6650 234.9450 155.6650 236.9450 ;
        RECT 162.1800 234.9450 164.1800 236.9450 ;
        RECT 170.6950 234.9450 172.6950 236.9450 ;
        RECT 145.1500 242.0400 147.1500 244.0400 ;
        RECT 153.6650 242.0400 155.6650 244.0400 ;
        RECT 162.1800 242.0400 164.1800 244.0400 ;
        RECT 170.6950 242.0400 172.6950 244.0400 ;
        RECT 204.7550 220.7550 206.7550 222.7550 ;
        RECT 196.2400 220.7550 198.2400 222.7550 ;
        RECT 187.7250 220.7550 189.7250 222.7550 ;
        RECT 179.2100 220.7550 181.2100 222.7550 ;
        RECT 204.7550 213.6600 206.7550 215.6600 ;
        RECT 196.2400 213.6600 198.2400 215.6600 ;
        RECT 187.7250 213.6600 189.7250 215.6600 ;
        RECT 179.2100 213.6600 181.2100 215.6600 ;
        RECT 187.7250 227.8500 189.7250 229.8500 ;
        RECT 179.2100 227.8500 181.2100 229.8500 ;
        RECT 196.2400 227.8500 198.2400 229.8500 ;
        RECT 204.7550 227.8500 206.7550 229.8500 ;
        RECT 179.2100 234.9450 181.2100 236.9450 ;
        RECT 187.7250 234.9450 189.7250 236.9450 ;
        RECT 196.2400 234.9450 198.2400 236.9450 ;
        RECT 204.7550 234.9450 206.7550 236.9450 ;
        RECT 179.2100 242.0400 181.2100 244.0400 ;
        RECT 187.7250 242.0400 189.7250 244.0400 ;
        RECT 196.2400 242.0400 198.2400 244.0400 ;
        RECT 204.7550 242.0400 206.7550 244.0400 ;
        RECT 170.6950 256.2300 172.6950 258.2300 ;
        RECT 162.1800 256.2300 164.1800 258.2300 ;
        RECT 153.6650 256.2300 155.6650 258.2300 ;
        RECT 145.1500 256.2300 147.1500 258.2300 ;
        RECT 170.6950 249.1350 172.6950 251.1350 ;
        RECT 162.1800 249.1350 164.1800 251.1350 ;
        RECT 153.6650 249.1350 155.6650 251.1350 ;
        RECT 145.1500 249.1350 147.1500 251.1350 ;
        RECT 153.6650 263.3250 155.6650 265.3250 ;
        RECT 145.1500 263.3250 147.1500 265.3250 ;
        RECT 162.1800 263.3250 164.1800 265.3250 ;
        RECT 170.6950 263.3250 172.6950 265.3250 ;
        RECT 145.1500 270.4200 147.1500 272.4200 ;
        RECT 153.6650 270.4200 155.6650 272.4200 ;
        RECT 162.1800 270.4200 164.1800 272.4200 ;
        RECT 170.6950 270.4200 172.6950 272.4200 ;
        RECT 145.1500 277.5150 147.1500 279.5150 ;
        RECT 153.6650 277.5150 155.6650 279.5150 ;
        RECT 162.1800 277.5150 164.1800 279.5150 ;
        RECT 170.6950 277.5150 172.6950 279.5150 ;
        RECT 204.7550 256.2300 206.7550 258.2300 ;
        RECT 196.2400 256.2300 198.2400 258.2300 ;
        RECT 187.7250 256.2300 189.7250 258.2300 ;
        RECT 179.2100 256.2300 181.2100 258.2300 ;
        RECT 204.7550 249.1350 206.7550 251.1350 ;
        RECT 196.2400 249.1350 198.2400 251.1350 ;
        RECT 187.7250 249.1350 189.7250 251.1350 ;
        RECT 179.2100 249.1350 181.2100 251.1350 ;
        RECT 187.7250 263.3250 189.7250 265.3250 ;
        RECT 179.2100 263.3250 181.2100 265.3250 ;
        RECT 196.2400 263.3250 198.2400 265.3250 ;
        RECT 204.7550 263.3250 206.7550 265.3250 ;
        RECT 179.2100 270.4200 181.2100 272.4200 ;
        RECT 187.7250 270.4200 189.7250 272.4200 ;
        RECT 196.2400 270.4200 198.2400 272.4200 ;
        RECT 204.7550 270.4200 206.7550 272.4200 ;
        RECT 179.2100 277.5150 181.2100 279.5150 ;
        RECT 187.7250 277.5150 189.7250 279.5150 ;
        RECT 196.2400 277.5150 198.2400 279.5150 ;
        RECT 204.7550 277.5150 206.7550 279.5150 ;
        RECT 238.8150 220.7550 240.8150 222.7550 ;
        RECT 230.3000 220.7550 232.3000 222.7550 ;
        RECT 221.7850 220.7550 223.7850 222.7550 ;
        RECT 213.2700 220.7550 215.2700 222.7550 ;
        RECT 238.8150 213.6600 240.8150 215.6600 ;
        RECT 230.3000 213.6600 232.3000 215.6600 ;
        RECT 221.7850 213.6600 223.7850 215.6600 ;
        RECT 213.2700 213.6600 215.2700 215.6600 ;
        RECT 221.7850 227.8500 223.7850 229.8500 ;
        RECT 213.2700 227.8500 215.2700 229.8500 ;
        RECT 230.3000 227.8500 232.3000 229.8500 ;
        RECT 238.8150 227.8500 240.8150 229.8500 ;
        RECT 213.2700 234.9450 215.2700 236.9450 ;
        RECT 221.7850 234.9450 223.7850 236.9450 ;
        RECT 230.3000 234.9450 232.3000 236.9450 ;
        RECT 238.8150 234.9450 240.8150 236.9450 ;
        RECT 213.2700 242.0400 215.2700 244.0400 ;
        RECT 221.7850 242.0400 223.7850 244.0400 ;
        RECT 230.3000 242.0400 232.3000 244.0400 ;
        RECT 238.8150 242.0400 240.8150 244.0400 ;
        RECT 272.8750 220.7550 274.8750 222.7550 ;
        RECT 264.3600 220.7550 266.3600 222.7550 ;
        RECT 255.8450 220.7550 257.8450 222.7550 ;
        RECT 247.3300 220.7550 249.3300 222.7550 ;
        RECT 272.8750 213.6600 274.8750 215.6600 ;
        RECT 264.3600 213.6600 266.3600 215.6600 ;
        RECT 255.8450 213.6600 257.8450 215.6600 ;
        RECT 247.3300 213.6600 249.3300 215.6600 ;
        RECT 255.8450 227.8500 257.8450 229.8500 ;
        RECT 247.3300 227.8500 249.3300 229.8500 ;
        RECT 264.3600 227.8500 266.3600 229.8500 ;
        RECT 272.8750 227.8500 274.8750 229.8500 ;
        RECT 247.3300 234.9450 249.3300 236.9450 ;
        RECT 255.8450 234.9450 257.8450 236.9450 ;
        RECT 264.3600 234.9450 266.3600 236.9450 ;
        RECT 272.8750 234.9450 274.8750 236.9450 ;
        RECT 247.3300 242.0400 249.3300 244.0400 ;
        RECT 255.8450 242.0400 257.8450 244.0400 ;
        RECT 264.3600 242.0400 266.3600 244.0400 ;
        RECT 272.8750 242.0400 274.8750 244.0400 ;
        RECT 238.8150 256.2300 240.8150 258.2300 ;
        RECT 230.3000 256.2300 232.3000 258.2300 ;
        RECT 221.7850 256.2300 223.7850 258.2300 ;
        RECT 213.2700 256.2300 215.2700 258.2300 ;
        RECT 238.8150 249.1350 240.8150 251.1350 ;
        RECT 230.3000 249.1350 232.3000 251.1350 ;
        RECT 221.7850 249.1350 223.7850 251.1350 ;
        RECT 213.2700 249.1350 215.2700 251.1350 ;
        RECT 221.7850 263.3250 223.7850 265.3250 ;
        RECT 213.2700 263.3250 215.2700 265.3250 ;
        RECT 230.3000 263.3250 232.3000 265.3250 ;
        RECT 238.8150 263.3250 240.8150 265.3250 ;
        RECT 213.2700 270.4200 215.2700 272.4200 ;
        RECT 221.7850 270.4200 223.7850 272.4200 ;
        RECT 230.3000 270.4200 232.3000 272.4200 ;
        RECT 238.8150 270.4200 240.8150 272.4200 ;
        RECT 213.2700 277.5150 215.2700 279.5150 ;
        RECT 221.7850 277.5150 223.7850 279.5150 ;
        RECT 230.3000 277.5150 232.3000 279.5150 ;
        RECT 238.8150 277.5150 240.8150 279.5150 ;
        RECT 272.8750 256.2300 274.8750 258.2300 ;
        RECT 264.3600 256.2300 266.3600 258.2300 ;
        RECT 255.8450 256.2300 257.8450 258.2300 ;
        RECT 247.3300 256.2300 249.3300 258.2300 ;
        RECT 272.8750 249.1350 274.8750 251.1350 ;
        RECT 264.3600 249.1350 266.3600 251.1350 ;
        RECT 255.8450 249.1350 257.8450 251.1350 ;
        RECT 247.3300 249.1350 249.3300 251.1350 ;
        RECT 255.8450 263.3250 257.8450 265.3250 ;
        RECT 247.3300 263.3250 249.3300 265.3250 ;
        RECT 264.3600 263.3250 266.3600 265.3250 ;
        RECT 272.8750 263.3250 274.8750 265.3250 ;
        RECT 247.3300 270.4200 249.3300 272.4200 ;
        RECT 255.8450 270.4200 257.8450 272.4200 ;
        RECT 264.3600 270.4200 266.3600 272.4200 ;
        RECT 272.8750 270.4200 274.8750 272.4200 ;
        RECT 247.3300 277.5150 249.3300 279.5150 ;
        RECT 255.8450 277.5150 257.8450 279.5150 ;
        RECT 264.3600 277.5150 266.3600 279.5150 ;
        RECT 272.8750 277.5150 274.8750 279.5150 ;
        RECT 281.3900 64.6650 283.3900 66.6650 ;
        RECT 289.9050 64.6650 291.9050 66.6650 ;
        RECT 298.4200 64.6650 300.4200 66.6650 ;
        RECT 306.9350 64.6650 308.9350 66.6650 ;
        RECT 344.0000 44.0000 346.0000 45.3800 ;
        RECT 344.0000 50.4750 346.0000 52.4750 ;
        RECT 323.9650 64.6650 325.9650 66.6650 ;
        RECT 315.4500 64.6650 317.4500 66.6650 ;
        RECT 344.0000 64.6650 346.0000 66.6650 ;
        RECT 344.0000 57.5700 346.0000 59.5700 ;
        RECT 394.0000 50.4750 396.0000 52.4750 ;
        RECT 394.0000 44.0000 396.0000 45.3800 ;
        RECT 394.0000 64.6650 396.0000 66.6650 ;
        RECT 394.0000 57.5700 396.0000 59.5700 ;
        RECT 414.1500 64.6650 416.1500 66.6650 ;
        RECT 281.3900 85.9500 283.3900 87.9500 ;
        RECT 289.9050 85.9500 291.9050 87.9500 ;
        RECT 298.4200 85.9500 300.4200 87.9500 ;
        RECT 306.9350 85.9500 308.9350 87.9500 ;
        RECT 306.9350 78.8550 308.9350 80.8550 ;
        RECT 298.4200 78.8550 300.4200 80.8550 ;
        RECT 289.9050 78.8550 291.9050 80.8550 ;
        RECT 281.3900 78.8550 283.3900 80.8550 ;
        RECT 306.9350 71.7600 308.9350 73.7600 ;
        RECT 298.4200 71.7600 300.4200 73.7600 ;
        RECT 289.9050 71.7600 291.9050 73.7600 ;
        RECT 281.3900 71.7600 283.3900 73.7600 ;
        RECT 281.3900 93.0450 283.3900 95.0450 ;
        RECT 289.9050 93.0450 291.9050 95.0450 ;
        RECT 298.4200 93.0450 300.4200 95.0450 ;
        RECT 306.9350 93.0450 308.9350 95.0450 ;
        RECT 281.3900 100.1400 283.3900 102.1400 ;
        RECT 289.9050 100.1400 291.9050 102.1400 ;
        RECT 298.4200 100.1400 300.4200 102.1400 ;
        RECT 306.9350 100.1400 308.9350 102.1400 ;
        RECT 344.0000 85.9500 346.0000 87.9500 ;
        RECT 315.4500 85.9500 317.4500 87.9500 ;
        RECT 323.9650 85.9500 325.9650 87.9500 ;
        RECT 323.9650 78.8550 325.9650 80.8550 ;
        RECT 315.4500 78.8550 317.4500 80.8550 ;
        RECT 323.9650 71.7600 325.9650 73.7600 ;
        RECT 315.4500 71.7600 317.4500 73.7600 ;
        RECT 344.0000 78.8550 346.0000 80.8550 ;
        RECT 344.0000 71.7600 346.0000 73.7600 ;
        RECT 323.9650 100.1400 325.9650 102.1400 ;
        RECT 315.4500 100.1400 317.4500 102.1400 ;
        RECT 323.9650 93.0450 325.9650 95.0450 ;
        RECT 315.4500 93.0450 317.4500 95.0450 ;
        RECT 344.0000 100.1400 346.0000 102.1400 ;
        RECT 344.0000 93.0450 346.0000 95.0450 ;
        RECT 281.3900 121.4250 283.3900 123.4250 ;
        RECT 289.9050 121.4250 291.9050 123.4250 ;
        RECT 298.4200 121.4250 300.4200 123.4250 ;
        RECT 306.9350 121.4250 308.9350 123.4250 ;
        RECT 306.9350 114.3300 308.9350 116.3300 ;
        RECT 298.4200 114.3300 300.4200 116.3300 ;
        RECT 289.9050 114.3300 291.9050 116.3300 ;
        RECT 281.3900 114.3300 283.3900 116.3300 ;
        RECT 306.9350 107.2350 308.9350 109.2350 ;
        RECT 298.4200 107.2350 300.4200 109.2350 ;
        RECT 289.9050 107.2350 291.9050 109.2350 ;
        RECT 281.3900 107.2350 283.3900 109.2350 ;
        RECT 281.3900 128.5200 283.3900 130.5200 ;
        RECT 289.9050 128.5200 291.9050 130.5200 ;
        RECT 298.4200 128.5200 300.4200 130.5200 ;
        RECT 306.9350 128.5200 308.9350 130.5200 ;
        RECT 281.3900 135.6150 283.3900 137.6150 ;
        RECT 289.9050 135.6150 291.9050 137.6150 ;
        RECT 298.4200 135.6150 300.4200 137.6150 ;
        RECT 306.9350 135.6150 308.9350 137.6150 ;
        RECT 344.0000 121.4250 346.0000 123.4250 ;
        RECT 315.4500 121.4250 317.4500 123.4250 ;
        RECT 323.9650 121.4250 325.9650 123.4250 ;
        RECT 323.9650 114.3300 325.9650 116.3300 ;
        RECT 315.4500 114.3300 317.4500 116.3300 ;
        RECT 323.9650 107.2350 325.9650 109.2350 ;
        RECT 315.4500 107.2350 317.4500 109.2350 ;
        RECT 344.0000 107.2350 346.0000 109.2350 ;
        RECT 344.0000 114.3300 346.0000 116.3300 ;
        RECT 323.9650 128.5200 325.9650 130.5200 ;
        RECT 315.4500 128.5200 317.4500 130.5200 ;
        RECT 315.4500 135.6150 317.4500 137.6150 ;
        RECT 323.9650 135.6150 325.9650 137.6150 ;
        RECT 344.0000 128.5200 346.0000 130.5200 ;
        RECT 344.0000 135.6150 346.0000 137.6150 ;
        RECT 394.0000 85.9500 396.0000 87.9500 ;
        RECT 414.1500 85.9500 416.1500 87.9500 ;
        RECT 394.0000 71.7600 396.0000 73.7600 ;
        RECT 394.0000 78.8550 396.0000 80.8550 ;
        RECT 414.1500 71.7600 416.1500 73.7600 ;
        RECT 414.1500 78.8550 416.1500 80.8550 ;
        RECT 394.0000 93.0450 396.0000 95.0450 ;
        RECT 394.0000 100.1400 396.0000 102.1400 ;
        RECT 414.1500 93.0450 416.1500 95.0450 ;
        RECT 414.1500 100.1400 416.1500 102.1400 ;
        RECT 394.0000 121.4250 396.0000 123.4250 ;
        RECT 414.1500 121.4250 416.1500 123.4250 ;
        RECT 394.0000 114.3300 396.0000 116.3300 ;
        RECT 394.0000 107.2350 396.0000 109.2350 ;
        RECT 414.1500 114.3300 416.1500 116.3300 ;
        RECT 414.1500 107.2350 416.1500 109.2350 ;
        RECT 394.0000 135.6150 396.0000 137.6150 ;
        RECT 394.0000 128.5200 396.0000 130.5200 ;
        RECT 414.1500 135.6150 416.1500 137.6150 ;
        RECT 414.1500 128.5200 416.1500 130.5200 ;
        RECT 487.5000 64.6650 489.5000 66.6650 ;
        RECT 479.3500 64.6650 481.3500 66.6650 ;
        RECT 471.2000 64.6650 473.2000 66.6650 ;
        RECT 463.0500 64.6650 465.0500 66.6650 ;
        RECT 454.9000 64.6650 456.9000 66.6650 ;
        RECT 446.7500 64.6650 448.7500 66.6650 ;
        RECT 438.6000 64.6650 440.6000 66.6650 ;
        RECT 430.4500 64.6650 432.4500 66.6650 ;
        RECT 422.3000 64.6650 424.3000 66.6650 ;
        RECT 520.1000 64.6650 522.1000 66.6650 ;
        RECT 511.9500 64.6650 513.9500 66.6650 ;
        RECT 503.8000 64.6650 505.8000 66.6650 ;
        RECT 495.6500 64.6650 497.6500 66.6650 ;
        RECT 528.2500 64.6650 530.2500 66.6650 ;
        RECT 536.4000 64.6650 538.4000 66.6650 ;
        RECT 544.5500 64.6650 546.5500 66.6650 ;
        RECT 552.7000 64.6650 554.7000 66.6650 ;
        RECT 454.9000 71.7600 456.9000 73.7600 ;
        RECT 454.9000 78.8550 456.9000 80.8550 ;
        RECT 454.9000 85.9500 456.9000 87.9500 ;
        RECT 454.9000 93.0450 456.9000 95.0450 ;
        RECT 454.9000 100.1400 456.9000 102.1400 ;
        RECT 422.3000 85.9500 424.3000 87.9500 ;
        RECT 430.4500 85.9500 432.4500 87.9500 ;
        RECT 438.6000 85.9500 440.6000 87.9500 ;
        RECT 446.7500 85.9500 448.7500 87.9500 ;
        RECT 446.7500 78.8550 448.7500 80.8550 ;
        RECT 438.6000 78.8550 440.6000 80.8550 ;
        RECT 430.4500 78.8550 432.4500 80.8550 ;
        RECT 422.3000 78.8550 424.3000 80.8550 ;
        RECT 446.7500 71.7600 448.7500 73.7600 ;
        RECT 438.6000 71.7600 440.6000 73.7600 ;
        RECT 430.4500 71.7600 432.4500 73.7600 ;
        RECT 422.3000 71.7600 424.3000 73.7600 ;
        RECT 422.3000 93.0450 424.3000 95.0450 ;
        RECT 430.4500 93.0450 432.4500 95.0450 ;
        RECT 438.6000 93.0450 440.6000 95.0450 ;
        RECT 446.7500 93.0450 448.7500 95.0450 ;
        RECT 422.3000 100.1400 424.3000 102.1400 ;
        RECT 430.4500 100.1400 432.4500 102.1400 ;
        RECT 438.6000 100.1400 440.6000 102.1400 ;
        RECT 446.7500 100.1400 448.7500 102.1400 ;
        RECT 463.0500 85.9500 465.0500 87.9500 ;
        RECT 471.2000 85.9500 473.2000 87.9500 ;
        RECT 479.3500 85.9500 481.3500 87.9500 ;
        RECT 487.5000 85.9500 489.5000 87.9500 ;
        RECT 487.5000 78.8550 489.5000 80.8550 ;
        RECT 479.3500 78.8550 481.3500 80.8550 ;
        RECT 471.2000 78.8550 473.2000 80.8550 ;
        RECT 463.0500 78.8550 465.0500 80.8550 ;
        RECT 487.5000 71.7600 489.5000 73.7600 ;
        RECT 479.3500 71.7600 481.3500 73.7600 ;
        RECT 471.2000 71.7600 473.2000 73.7600 ;
        RECT 463.0500 71.7600 465.0500 73.7600 ;
        RECT 463.0500 93.0450 465.0500 95.0450 ;
        RECT 471.2000 93.0450 473.2000 95.0450 ;
        RECT 479.3500 93.0450 481.3500 95.0450 ;
        RECT 487.5000 93.0450 489.5000 95.0450 ;
        RECT 463.0500 100.1400 465.0500 102.1400 ;
        RECT 471.2000 100.1400 473.2000 102.1400 ;
        RECT 479.3500 100.1400 481.3500 102.1400 ;
        RECT 487.5000 100.1400 489.5000 102.1400 ;
        RECT 454.9000 107.2350 456.9000 109.2350 ;
        RECT 454.9000 114.3300 456.9000 116.3300 ;
        RECT 454.9000 121.4250 456.9000 123.4250 ;
        RECT 454.9000 128.5200 456.9000 130.5200 ;
        RECT 454.9000 135.6150 456.9000 137.6150 ;
        RECT 422.3000 121.4250 424.3000 123.4250 ;
        RECT 430.4500 121.4250 432.4500 123.4250 ;
        RECT 438.6000 121.4250 440.6000 123.4250 ;
        RECT 446.7500 121.4250 448.7500 123.4250 ;
        RECT 446.7500 114.3300 448.7500 116.3300 ;
        RECT 438.6000 114.3300 440.6000 116.3300 ;
        RECT 430.4500 114.3300 432.4500 116.3300 ;
        RECT 422.3000 114.3300 424.3000 116.3300 ;
        RECT 446.7500 107.2350 448.7500 109.2350 ;
        RECT 438.6000 107.2350 440.6000 109.2350 ;
        RECT 430.4500 107.2350 432.4500 109.2350 ;
        RECT 422.3000 107.2350 424.3000 109.2350 ;
        RECT 422.3000 128.5200 424.3000 130.5200 ;
        RECT 430.4500 128.5200 432.4500 130.5200 ;
        RECT 438.6000 128.5200 440.6000 130.5200 ;
        RECT 446.7500 128.5200 448.7500 130.5200 ;
        RECT 422.3000 135.6150 424.3000 137.6150 ;
        RECT 430.4500 135.6150 432.4500 137.6150 ;
        RECT 438.6000 135.6150 440.6000 137.6150 ;
        RECT 446.7500 135.6150 448.7500 137.6150 ;
        RECT 463.0500 121.4250 465.0500 123.4250 ;
        RECT 471.2000 121.4250 473.2000 123.4250 ;
        RECT 479.3500 121.4250 481.3500 123.4250 ;
        RECT 487.5000 121.4250 489.5000 123.4250 ;
        RECT 487.5000 114.3300 489.5000 116.3300 ;
        RECT 479.3500 114.3300 481.3500 116.3300 ;
        RECT 471.2000 114.3300 473.2000 116.3300 ;
        RECT 463.0500 114.3300 465.0500 116.3300 ;
        RECT 487.5000 107.2350 489.5000 109.2350 ;
        RECT 479.3500 107.2350 481.3500 109.2350 ;
        RECT 471.2000 107.2350 473.2000 109.2350 ;
        RECT 463.0500 107.2350 465.0500 109.2350 ;
        RECT 463.0500 128.5200 465.0500 130.5200 ;
        RECT 471.2000 128.5200 473.2000 130.5200 ;
        RECT 479.3500 128.5200 481.3500 130.5200 ;
        RECT 487.5000 128.5200 489.5000 130.5200 ;
        RECT 463.0500 135.6150 465.0500 137.6150 ;
        RECT 471.2000 135.6150 473.2000 137.6150 ;
        RECT 479.3500 135.6150 481.3500 137.6150 ;
        RECT 487.5000 135.6150 489.5000 137.6150 ;
        RECT 495.6500 85.9500 497.6500 87.9500 ;
        RECT 503.8000 85.9500 505.8000 87.9500 ;
        RECT 511.9500 85.9500 513.9500 87.9500 ;
        RECT 520.1000 85.9500 522.1000 87.9500 ;
        RECT 520.1000 78.8550 522.1000 80.8550 ;
        RECT 511.9500 78.8550 513.9500 80.8550 ;
        RECT 503.8000 78.8550 505.8000 80.8550 ;
        RECT 495.6500 78.8550 497.6500 80.8550 ;
        RECT 520.1000 71.7600 522.1000 73.7600 ;
        RECT 511.9500 71.7600 513.9500 73.7600 ;
        RECT 503.8000 71.7600 505.8000 73.7600 ;
        RECT 495.6500 71.7600 497.6500 73.7600 ;
        RECT 495.6500 93.0450 497.6500 95.0450 ;
        RECT 503.8000 93.0450 505.8000 95.0450 ;
        RECT 511.9500 93.0450 513.9500 95.0450 ;
        RECT 520.1000 93.0450 522.1000 95.0450 ;
        RECT 495.6500 100.1400 497.6500 102.1400 ;
        RECT 503.8000 100.1400 505.8000 102.1400 ;
        RECT 511.9500 100.1400 513.9500 102.1400 ;
        RECT 520.1000 100.1400 522.1000 102.1400 ;
        RECT 528.2500 85.9500 530.2500 87.9500 ;
        RECT 536.4000 85.9500 538.4000 87.9500 ;
        RECT 544.5500 85.9500 546.5500 87.9500 ;
        RECT 552.7000 85.9500 554.7000 87.9500 ;
        RECT 552.7000 78.8550 554.7000 80.8550 ;
        RECT 544.5500 78.8550 546.5500 80.8550 ;
        RECT 536.4000 78.8550 538.4000 80.8550 ;
        RECT 528.2500 78.8550 530.2500 80.8550 ;
        RECT 552.7000 71.7600 554.7000 73.7600 ;
        RECT 544.5500 71.7600 546.5500 73.7600 ;
        RECT 536.4000 71.7600 538.4000 73.7600 ;
        RECT 528.2500 71.7600 530.2500 73.7600 ;
        RECT 528.2500 93.0450 530.2500 95.0450 ;
        RECT 536.4000 93.0450 538.4000 95.0450 ;
        RECT 544.5500 93.0450 546.5500 95.0450 ;
        RECT 552.7000 93.0450 554.7000 95.0450 ;
        RECT 528.2500 100.1400 530.2500 102.1400 ;
        RECT 536.4000 100.1400 538.4000 102.1400 ;
        RECT 544.5500 100.1400 546.5500 102.1400 ;
        RECT 552.7000 100.1400 554.7000 102.1400 ;
        RECT 495.6500 121.4250 497.6500 123.4250 ;
        RECT 503.8000 121.4250 505.8000 123.4250 ;
        RECT 511.9500 121.4250 513.9500 123.4250 ;
        RECT 520.1000 121.4250 522.1000 123.4250 ;
        RECT 520.1000 114.3300 522.1000 116.3300 ;
        RECT 511.9500 114.3300 513.9500 116.3300 ;
        RECT 503.8000 114.3300 505.8000 116.3300 ;
        RECT 495.6500 114.3300 497.6500 116.3300 ;
        RECT 520.1000 107.2350 522.1000 109.2350 ;
        RECT 511.9500 107.2350 513.9500 109.2350 ;
        RECT 503.8000 107.2350 505.8000 109.2350 ;
        RECT 495.6500 107.2350 497.6500 109.2350 ;
        RECT 495.6500 128.5200 497.6500 130.5200 ;
        RECT 503.8000 128.5200 505.8000 130.5200 ;
        RECT 511.9500 128.5200 513.9500 130.5200 ;
        RECT 520.1000 128.5200 522.1000 130.5200 ;
        RECT 495.6500 135.6150 497.6500 137.6150 ;
        RECT 503.8000 135.6150 505.8000 137.6150 ;
        RECT 511.9500 135.6150 513.9500 137.6150 ;
        RECT 520.1000 135.6150 522.1000 137.6150 ;
        RECT 528.2500 121.4250 530.2500 123.4250 ;
        RECT 536.4000 121.4250 538.4000 123.4250 ;
        RECT 544.5500 121.4250 546.5500 123.4250 ;
        RECT 552.7000 121.4250 554.7000 123.4250 ;
        RECT 552.7000 114.3300 554.7000 116.3300 ;
        RECT 544.5500 114.3300 546.5500 116.3300 ;
        RECT 536.4000 114.3300 538.4000 116.3300 ;
        RECT 528.2500 114.3300 530.2500 116.3300 ;
        RECT 552.7000 107.2350 554.7000 109.2350 ;
        RECT 544.5500 107.2350 546.5500 109.2350 ;
        RECT 536.4000 107.2350 538.4000 109.2350 ;
        RECT 528.2500 107.2350 530.2500 109.2350 ;
        RECT 528.2500 128.5200 530.2500 130.5200 ;
        RECT 536.4000 128.5200 538.4000 130.5200 ;
        RECT 544.5500 128.5200 546.5500 130.5200 ;
        RECT 552.7000 128.5200 554.7000 130.5200 ;
        RECT 528.2500 135.6150 530.2500 137.6150 ;
        RECT 536.4000 135.6150 538.4000 137.6150 ;
        RECT 544.5500 135.6150 546.5500 137.6150 ;
        RECT 552.7000 135.6150 554.7000 137.6150 ;
        RECT 281.3900 156.9000 283.3900 158.9000 ;
        RECT 289.9050 156.9000 291.9050 158.9000 ;
        RECT 298.4200 156.9000 300.4200 158.9000 ;
        RECT 306.9350 156.9000 308.9350 158.9000 ;
        RECT 306.9350 149.8050 308.9350 151.8050 ;
        RECT 298.4200 149.8050 300.4200 151.8050 ;
        RECT 289.9050 149.8050 291.9050 151.8050 ;
        RECT 281.3900 149.8050 283.3900 151.8050 ;
        RECT 306.9350 142.7100 308.9350 144.7100 ;
        RECT 298.4200 142.7100 300.4200 144.7100 ;
        RECT 289.9050 142.7100 291.9050 144.7100 ;
        RECT 281.3900 142.7100 283.3900 144.7100 ;
        RECT 281.3900 163.9950 283.3900 165.9950 ;
        RECT 289.9050 163.9950 291.9050 165.9950 ;
        RECT 298.4200 163.9950 300.4200 165.9950 ;
        RECT 306.9350 163.9950 308.9350 165.9950 ;
        RECT 281.3900 171.0900 283.3900 173.0900 ;
        RECT 289.9050 171.0900 291.9050 173.0900 ;
        RECT 298.4200 171.0900 300.4200 173.0900 ;
        RECT 306.9350 171.0900 308.9350 173.0900 ;
        RECT 344.0000 156.9000 346.0000 158.9000 ;
        RECT 315.4500 156.9000 317.4500 158.9000 ;
        RECT 323.9650 156.9000 325.9650 158.9000 ;
        RECT 323.9650 149.8050 325.9650 151.8050 ;
        RECT 315.4500 149.8050 317.4500 151.8050 ;
        RECT 323.9650 142.7100 325.9650 144.7100 ;
        RECT 315.4500 142.7100 317.4500 144.7100 ;
        RECT 344.0000 142.7100 346.0000 144.7100 ;
        RECT 344.0000 149.8050 346.0000 151.8050 ;
        RECT 323.9650 171.0900 325.9650 173.0900 ;
        RECT 315.4500 171.0900 317.4500 173.0900 ;
        RECT 323.9650 163.9950 325.9650 165.9950 ;
        RECT 315.4500 163.9950 317.4500 165.9950 ;
        RECT 344.0000 163.9950 346.0000 165.9950 ;
        RECT 344.0000 171.0900 346.0000 173.0900 ;
        RECT 281.3900 192.3750 283.3900 194.3750 ;
        RECT 289.9050 192.3750 291.9050 194.3750 ;
        RECT 298.4200 192.3750 300.4200 194.3750 ;
        RECT 306.9350 192.3750 308.9350 194.3750 ;
        RECT 306.9350 185.2800 308.9350 187.2800 ;
        RECT 298.4200 185.2800 300.4200 187.2800 ;
        RECT 289.9050 185.2800 291.9050 187.2800 ;
        RECT 281.3900 185.2800 283.3900 187.2800 ;
        RECT 306.9350 178.1850 308.9350 180.1850 ;
        RECT 298.4200 178.1850 300.4200 180.1850 ;
        RECT 289.9050 178.1850 291.9050 180.1850 ;
        RECT 281.3900 178.1850 283.3900 180.1850 ;
        RECT 281.3900 199.4700 283.3900 201.4700 ;
        RECT 289.9050 199.4700 291.9050 201.4700 ;
        RECT 298.4200 199.4700 300.4200 201.4700 ;
        RECT 306.9350 199.4700 308.9350 201.4700 ;
        RECT 281.3900 206.5650 283.3900 208.5650 ;
        RECT 289.9050 206.5650 291.9050 208.5650 ;
        RECT 298.4200 206.5650 300.4200 208.5650 ;
        RECT 306.9350 206.5650 308.9350 208.5650 ;
        RECT 344.0000 192.3750 346.0000 194.3750 ;
        RECT 315.4500 192.3750 317.4500 194.3750 ;
        RECT 323.9650 192.3750 325.9650 194.3750 ;
        RECT 315.4500 185.2800 317.4500 187.2800 ;
        RECT 323.9650 178.1850 325.9650 180.1850 ;
        RECT 315.4500 178.1850 317.4500 180.1850 ;
        RECT 323.9650 185.2800 325.9650 187.2800 ;
        RECT 344.0000 178.1850 346.0000 180.1850 ;
        RECT 344.0000 185.2800 346.0000 187.2800 ;
        RECT 323.9650 199.4700 325.9650 201.4700 ;
        RECT 315.4500 199.4700 317.4500 201.4700 ;
        RECT 315.4500 206.5650 317.4500 208.5650 ;
        RECT 323.9650 206.5650 325.9650 208.5650 ;
        RECT 344.0000 199.4700 346.0000 201.4700 ;
        RECT 344.0000 206.5650 346.0000 208.5650 ;
        RECT 394.0000 156.9000 396.0000 158.9000 ;
        RECT 414.1500 156.9000 416.1500 158.9000 ;
        RECT 394.0000 142.7100 396.0000 144.7100 ;
        RECT 394.0000 149.8050 396.0000 151.8050 ;
        RECT 414.1500 142.7100 416.1500 144.7100 ;
        RECT 414.1500 149.8050 416.1500 151.8050 ;
        RECT 394.0000 163.9950 396.0000 165.9950 ;
        RECT 394.0000 171.0900 396.0000 173.0900 ;
        RECT 414.1500 163.9950 416.1500 165.9950 ;
        RECT 414.1500 171.0900 416.1500 173.0900 ;
        RECT 394.0000 192.3750 396.0000 194.3750 ;
        RECT 414.1500 192.3750 416.1500 194.3750 ;
        RECT 394.0000 185.2800 396.0000 187.2800 ;
        RECT 394.0000 178.1850 396.0000 180.1850 ;
        RECT 414.1500 185.2800 416.1500 187.2800 ;
        RECT 414.1500 178.1850 416.1500 180.1850 ;
        RECT 394.0000 206.5650 396.0000 208.5650 ;
        RECT 394.0000 199.4700 396.0000 201.4700 ;
        RECT 414.1500 206.5650 416.1500 208.5650 ;
        RECT 414.1500 199.4700 416.1500 201.4700 ;
        RECT 306.9350 220.7550 308.9350 222.7550 ;
        RECT 298.4200 220.7550 300.4200 222.7550 ;
        RECT 289.9050 220.7550 291.9050 222.7550 ;
        RECT 281.3900 220.7550 283.3900 222.7550 ;
        RECT 306.9350 213.6600 308.9350 215.6600 ;
        RECT 298.4200 213.6600 300.4200 215.6600 ;
        RECT 289.9050 213.6600 291.9050 215.6600 ;
        RECT 281.3900 213.6600 283.3900 215.6600 ;
        RECT 289.9050 227.8500 291.9050 229.8500 ;
        RECT 281.3900 227.8500 283.3900 229.8500 ;
        RECT 298.4200 227.8500 300.4200 229.8500 ;
        RECT 306.9350 227.8500 308.9350 229.8500 ;
        RECT 281.3900 234.9450 283.3900 236.9450 ;
        RECT 289.9050 234.9450 291.9050 236.9450 ;
        RECT 298.4200 234.9450 300.4200 236.9450 ;
        RECT 306.9350 234.9450 308.9350 236.9450 ;
        RECT 281.3900 242.0400 283.3900 244.0400 ;
        RECT 289.9050 242.0400 291.9050 244.0400 ;
        RECT 298.4200 242.0400 300.4200 244.0400 ;
        RECT 306.9350 242.0400 308.9350 244.0400 ;
        RECT 323.9650 220.7550 325.9650 222.7550 ;
        RECT 315.4500 220.7550 317.4500 222.7550 ;
        RECT 323.9650 213.6600 325.9650 215.6600 ;
        RECT 315.4500 213.6600 317.4500 215.6600 ;
        RECT 344.0000 213.6600 346.0000 215.6600 ;
        RECT 344.0000 220.7550 346.0000 222.7550 ;
        RECT 315.4500 227.8500 317.4500 229.8500 ;
        RECT 323.9650 227.8500 325.9650 229.8500 ;
        RECT 315.4500 234.9450 317.4500 236.9450 ;
        RECT 323.9650 234.9450 325.9650 236.9450 ;
        RECT 315.4500 242.0400 317.4500 244.0400 ;
        RECT 323.9650 242.0400 325.9650 244.0400 ;
        RECT 344.0000 227.8500 346.0000 229.8500 ;
        RECT 344.0000 234.9450 346.0000 236.9450 ;
        RECT 344.0000 242.0400 346.0000 244.0400 ;
        RECT 306.9350 256.2300 308.9350 258.2300 ;
        RECT 298.4200 256.2300 300.4200 258.2300 ;
        RECT 289.9050 256.2300 291.9050 258.2300 ;
        RECT 281.3900 256.2300 283.3900 258.2300 ;
        RECT 306.9350 249.1350 308.9350 251.1350 ;
        RECT 298.4200 249.1350 300.4200 251.1350 ;
        RECT 289.9050 249.1350 291.9050 251.1350 ;
        RECT 281.3900 249.1350 283.3900 251.1350 ;
        RECT 289.9050 263.3250 291.9050 265.3250 ;
        RECT 281.3900 263.3250 283.3900 265.3250 ;
        RECT 298.4200 263.3250 300.4200 265.3250 ;
        RECT 306.9350 263.3250 308.9350 265.3250 ;
        RECT 281.3900 270.4200 283.3900 272.4200 ;
        RECT 289.9050 270.4200 291.9050 272.4200 ;
        RECT 298.4200 270.4200 300.4200 272.4200 ;
        RECT 306.9350 270.4200 308.9350 272.4200 ;
        RECT 281.3900 277.5150 283.3900 279.5150 ;
        RECT 289.9050 277.5150 291.9050 279.5150 ;
        RECT 298.4200 277.5150 300.4200 279.5150 ;
        RECT 306.9350 277.5150 308.9350 279.5150 ;
        RECT 323.9650 256.2300 325.9650 258.2300 ;
        RECT 315.4500 256.2300 317.4500 258.2300 ;
        RECT 323.9650 249.1350 325.9650 251.1350 ;
        RECT 315.4500 249.1350 317.4500 251.1350 ;
        RECT 344.0000 249.1350 346.0000 251.1350 ;
        RECT 344.0000 256.2300 346.0000 258.2300 ;
        RECT 323.9650 263.3250 325.9650 265.3250 ;
        RECT 315.4500 263.3250 317.4500 265.3250 ;
        RECT 315.4500 270.4200 317.4500 272.4200 ;
        RECT 323.9650 270.4200 325.9650 272.4200 ;
        RECT 315.4500 277.5150 317.4500 279.5150 ;
        RECT 323.9650 277.5150 325.9650 279.5150 ;
        RECT 344.0000 263.3250 346.0000 265.3250 ;
        RECT 344.0000 270.4200 346.0000 272.4200 ;
        RECT 344.0000 277.5150 346.0000 279.5150 ;
        RECT 394.0000 213.6600 396.0000 215.6600 ;
        RECT 394.0000 220.7550 396.0000 222.7550 ;
        RECT 414.1500 213.6600 416.1500 215.6600 ;
        RECT 414.1500 220.7550 416.1500 222.7550 ;
        RECT 394.0000 242.0400 396.0000 244.0400 ;
        RECT 394.0000 234.9450 396.0000 236.9450 ;
        RECT 394.0000 227.8500 396.0000 229.8500 ;
        RECT 414.1500 227.8500 416.1500 229.8500 ;
        RECT 414.1500 234.9450 416.1500 236.9450 ;
        RECT 414.1500 242.0400 416.1500 244.0400 ;
        RECT 394.0000 256.2300 396.0000 258.2300 ;
        RECT 394.0000 249.1350 396.0000 251.1350 ;
        RECT 414.1500 256.2300 416.1500 258.2300 ;
        RECT 414.1500 249.1350 416.1500 251.1350 ;
        RECT 394.0000 277.5150 396.0000 279.5150 ;
        RECT 394.0000 270.4200 396.0000 272.4200 ;
        RECT 394.0000 263.3250 396.0000 265.3250 ;
        RECT 414.1500 270.4200 416.1500 272.4200 ;
        RECT 414.1500 263.3250 416.1500 265.3250 ;
        RECT 414.1500 277.5150 416.1500 279.5150 ;
        RECT 454.9000 142.7100 456.9000 144.7100 ;
        RECT 454.9000 149.8050 456.9000 151.8050 ;
        RECT 454.9000 156.9000 456.9000 158.9000 ;
        RECT 454.9000 163.9950 456.9000 165.9950 ;
        RECT 454.9000 171.0900 456.9000 173.0900 ;
        RECT 422.3000 156.9000 424.3000 158.9000 ;
        RECT 430.4500 156.9000 432.4500 158.9000 ;
        RECT 438.6000 156.9000 440.6000 158.9000 ;
        RECT 446.7500 156.9000 448.7500 158.9000 ;
        RECT 446.7500 149.8050 448.7500 151.8050 ;
        RECT 438.6000 149.8050 440.6000 151.8050 ;
        RECT 430.4500 149.8050 432.4500 151.8050 ;
        RECT 422.3000 149.8050 424.3000 151.8050 ;
        RECT 446.7500 142.7100 448.7500 144.7100 ;
        RECT 438.6000 142.7100 440.6000 144.7100 ;
        RECT 430.4500 142.7100 432.4500 144.7100 ;
        RECT 422.3000 142.7100 424.3000 144.7100 ;
        RECT 422.3000 163.9950 424.3000 165.9950 ;
        RECT 430.4500 163.9950 432.4500 165.9950 ;
        RECT 438.6000 163.9950 440.6000 165.9950 ;
        RECT 446.7500 163.9950 448.7500 165.9950 ;
        RECT 422.3000 171.0900 424.3000 173.0900 ;
        RECT 430.4500 171.0900 432.4500 173.0900 ;
        RECT 438.6000 171.0900 440.6000 173.0900 ;
        RECT 446.7500 171.0900 448.7500 173.0900 ;
        RECT 463.0500 156.9000 465.0500 158.9000 ;
        RECT 471.2000 156.9000 473.2000 158.9000 ;
        RECT 479.3500 156.9000 481.3500 158.9000 ;
        RECT 487.5000 156.9000 489.5000 158.9000 ;
        RECT 487.5000 149.8050 489.5000 151.8050 ;
        RECT 479.3500 149.8050 481.3500 151.8050 ;
        RECT 471.2000 149.8050 473.2000 151.8050 ;
        RECT 463.0500 149.8050 465.0500 151.8050 ;
        RECT 487.5000 142.7100 489.5000 144.7100 ;
        RECT 479.3500 142.7100 481.3500 144.7100 ;
        RECT 471.2000 142.7100 473.2000 144.7100 ;
        RECT 463.0500 142.7100 465.0500 144.7100 ;
        RECT 463.0500 163.9950 465.0500 165.9950 ;
        RECT 471.2000 163.9950 473.2000 165.9950 ;
        RECT 479.3500 163.9950 481.3500 165.9950 ;
        RECT 487.5000 163.9950 489.5000 165.9950 ;
        RECT 463.0500 171.0900 465.0500 173.0900 ;
        RECT 471.2000 171.0900 473.2000 173.0900 ;
        RECT 479.3500 171.0900 481.3500 173.0900 ;
        RECT 487.5000 171.0900 489.5000 173.0900 ;
        RECT 454.9000 178.1850 456.9000 180.1850 ;
        RECT 454.9000 185.2800 456.9000 187.2800 ;
        RECT 454.9000 192.3750 456.9000 194.3750 ;
        RECT 454.9000 199.4700 456.9000 201.4700 ;
        RECT 454.9000 206.5650 456.9000 208.5650 ;
        RECT 422.3000 192.3750 424.3000 194.3750 ;
        RECT 430.4500 192.3750 432.4500 194.3750 ;
        RECT 438.6000 192.3750 440.6000 194.3750 ;
        RECT 446.7500 192.3750 448.7500 194.3750 ;
        RECT 446.7500 185.2800 448.7500 187.2800 ;
        RECT 438.6000 185.2800 440.6000 187.2800 ;
        RECT 430.4500 185.2800 432.4500 187.2800 ;
        RECT 422.3000 185.2800 424.3000 187.2800 ;
        RECT 446.7500 178.1850 448.7500 180.1850 ;
        RECT 438.6000 178.1850 440.6000 180.1850 ;
        RECT 430.4500 178.1850 432.4500 180.1850 ;
        RECT 422.3000 178.1850 424.3000 180.1850 ;
        RECT 422.3000 199.4700 424.3000 201.4700 ;
        RECT 430.4500 199.4700 432.4500 201.4700 ;
        RECT 438.6000 199.4700 440.6000 201.4700 ;
        RECT 446.7500 199.4700 448.7500 201.4700 ;
        RECT 422.3000 206.5650 424.3000 208.5650 ;
        RECT 430.4500 206.5650 432.4500 208.5650 ;
        RECT 438.6000 206.5650 440.6000 208.5650 ;
        RECT 446.7500 206.5650 448.7500 208.5650 ;
        RECT 463.0500 192.3750 465.0500 194.3750 ;
        RECT 471.2000 192.3750 473.2000 194.3750 ;
        RECT 479.3500 192.3750 481.3500 194.3750 ;
        RECT 487.5000 192.3750 489.5000 194.3750 ;
        RECT 487.5000 185.2800 489.5000 187.2800 ;
        RECT 479.3500 185.2800 481.3500 187.2800 ;
        RECT 471.2000 185.2800 473.2000 187.2800 ;
        RECT 463.0500 185.2800 465.0500 187.2800 ;
        RECT 487.5000 178.1850 489.5000 180.1850 ;
        RECT 479.3500 178.1850 481.3500 180.1850 ;
        RECT 471.2000 178.1850 473.2000 180.1850 ;
        RECT 463.0500 178.1850 465.0500 180.1850 ;
        RECT 463.0500 199.4700 465.0500 201.4700 ;
        RECT 471.2000 199.4700 473.2000 201.4700 ;
        RECT 479.3500 199.4700 481.3500 201.4700 ;
        RECT 487.5000 199.4700 489.5000 201.4700 ;
        RECT 463.0500 206.5650 465.0500 208.5650 ;
        RECT 471.2000 206.5650 473.2000 208.5650 ;
        RECT 479.3500 206.5650 481.3500 208.5650 ;
        RECT 487.5000 206.5650 489.5000 208.5650 ;
        RECT 495.6500 156.9000 497.6500 158.9000 ;
        RECT 503.8000 156.9000 505.8000 158.9000 ;
        RECT 511.9500 156.9000 513.9500 158.9000 ;
        RECT 520.1000 156.9000 522.1000 158.9000 ;
        RECT 520.1000 149.8050 522.1000 151.8050 ;
        RECT 511.9500 149.8050 513.9500 151.8050 ;
        RECT 503.8000 149.8050 505.8000 151.8050 ;
        RECT 495.6500 149.8050 497.6500 151.8050 ;
        RECT 520.1000 142.7100 522.1000 144.7100 ;
        RECT 511.9500 142.7100 513.9500 144.7100 ;
        RECT 503.8000 142.7100 505.8000 144.7100 ;
        RECT 495.6500 142.7100 497.6500 144.7100 ;
        RECT 495.6500 163.9950 497.6500 165.9950 ;
        RECT 503.8000 163.9950 505.8000 165.9950 ;
        RECT 511.9500 163.9950 513.9500 165.9950 ;
        RECT 520.1000 163.9950 522.1000 165.9950 ;
        RECT 495.6500 171.0900 497.6500 173.0900 ;
        RECT 503.8000 171.0900 505.8000 173.0900 ;
        RECT 511.9500 171.0900 513.9500 173.0900 ;
        RECT 520.1000 171.0900 522.1000 173.0900 ;
        RECT 528.2500 156.9000 530.2500 158.9000 ;
        RECT 536.4000 156.9000 538.4000 158.9000 ;
        RECT 544.5500 156.9000 546.5500 158.9000 ;
        RECT 552.7000 156.9000 554.7000 158.9000 ;
        RECT 552.7000 149.8050 554.7000 151.8050 ;
        RECT 544.5500 149.8050 546.5500 151.8050 ;
        RECT 536.4000 149.8050 538.4000 151.8050 ;
        RECT 528.2500 149.8050 530.2500 151.8050 ;
        RECT 552.7000 142.7100 554.7000 144.7100 ;
        RECT 544.5500 142.7100 546.5500 144.7100 ;
        RECT 536.4000 142.7100 538.4000 144.7100 ;
        RECT 528.2500 142.7100 530.2500 144.7100 ;
        RECT 528.2500 163.9950 530.2500 165.9950 ;
        RECT 536.4000 163.9950 538.4000 165.9950 ;
        RECT 544.5500 163.9950 546.5500 165.9950 ;
        RECT 552.7000 163.9950 554.7000 165.9950 ;
        RECT 528.2500 171.0900 530.2500 173.0900 ;
        RECT 536.4000 171.0900 538.4000 173.0900 ;
        RECT 544.5500 171.0900 546.5500 173.0900 ;
        RECT 552.7000 171.0900 554.7000 173.0900 ;
        RECT 495.6500 192.3750 497.6500 194.3750 ;
        RECT 503.8000 192.3750 505.8000 194.3750 ;
        RECT 511.9500 192.3750 513.9500 194.3750 ;
        RECT 520.1000 192.3750 522.1000 194.3750 ;
        RECT 520.1000 185.2800 522.1000 187.2800 ;
        RECT 511.9500 185.2800 513.9500 187.2800 ;
        RECT 503.8000 185.2800 505.8000 187.2800 ;
        RECT 495.6500 185.2800 497.6500 187.2800 ;
        RECT 520.1000 178.1850 522.1000 180.1850 ;
        RECT 511.9500 178.1850 513.9500 180.1850 ;
        RECT 503.8000 178.1850 505.8000 180.1850 ;
        RECT 495.6500 178.1850 497.6500 180.1850 ;
        RECT 495.6500 199.4700 497.6500 201.4700 ;
        RECT 503.8000 199.4700 505.8000 201.4700 ;
        RECT 511.9500 199.4700 513.9500 201.4700 ;
        RECT 520.1000 199.4700 522.1000 201.4700 ;
        RECT 495.6500 206.5650 497.6500 208.5650 ;
        RECT 503.8000 206.5650 505.8000 208.5650 ;
        RECT 511.9500 206.5650 513.9500 208.5650 ;
        RECT 520.1000 206.5650 522.1000 208.5650 ;
        RECT 528.2500 192.3750 530.2500 194.3750 ;
        RECT 536.4000 192.3750 538.4000 194.3750 ;
        RECT 544.5500 192.3750 546.5500 194.3750 ;
        RECT 552.7000 192.3750 554.7000 194.3750 ;
        RECT 552.7000 185.2800 554.7000 187.2800 ;
        RECT 544.5500 185.2800 546.5500 187.2800 ;
        RECT 536.4000 185.2800 538.4000 187.2800 ;
        RECT 528.2500 185.2800 530.2500 187.2800 ;
        RECT 552.7000 178.1850 554.7000 180.1850 ;
        RECT 544.5500 178.1850 546.5500 180.1850 ;
        RECT 536.4000 178.1850 538.4000 180.1850 ;
        RECT 528.2500 178.1850 530.2500 180.1850 ;
        RECT 528.2500 199.4700 530.2500 201.4700 ;
        RECT 536.4000 199.4700 538.4000 201.4700 ;
        RECT 544.5500 199.4700 546.5500 201.4700 ;
        RECT 552.7000 199.4700 554.7000 201.4700 ;
        RECT 528.2500 206.5650 530.2500 208.5650 ;
        RECT 536.4000 206.5650 538.4000 208.5650 ;
        RECT 544.5500 206.5650 546.5500 208.5650 ;
        RECT 552.7000 206.5650 554.7000 208.5650 ;
        RECT 454.9000 213.6600 456.9000 215.6600 ;
        RECT 454.9000 220.7550 456.9000 222.7550 ;
        RECT 454.9000 227.8500 456.9000 229.8500 ;
        RECT 454.9000 234.9450 456.9000 236.9450 ;
        RECT 454.9000 242.0400 456.9000 244.0400 ;
        RECT 446.7500 220.7550 448.7500 222.7550 ;
        RECT 438.6000 220.7550 440.6000 222.7550 ;
        RECT 430.4500 220.7550 432.4500 222.7550 ;
        RECT 422.3000 220.7550 424.3000 222.7550 ;
        RECT 446.7500 213.6600 448.7500 215.6600 ;
        RECT 438.6000 213.6600 440.6000 215.6600 ;
        RECT 430.4500 213.6600 432.4500 215.6600 ;
        RECT 422.3000 213.6600 424.3000 215.6600 ;
        RECT 430.4500 227.8500 432.4500 229.8500 ;
        RECT 422.3000 227.8500 424.3000 229.8500 ;
        RECT 438.6000 227.8500 440.6000 229.8500 ;
        RECT 446.7500 227.8500 448.7500 229.8500 ;
        RECT 422.3000 234.9450 424.3000 236.9450 ;
        RECT 430.4500 234.9450 432.4500 236.9450 ;
        RECT 438.6000 234.9450 440.6000 236.9450 ;
        RECT 446.7500 234.9450 448.7500 236.9450 ;
        RECT 422.3000 242.0400 424.3000 244.0400 ;
        RECT 430.4500 242.0400 432.4500 244.0400 ;
        RECT 438.6000 242.0400 440.6000 244.0400 ;
        RECT 446.7500 242.0400 448.7500 244.0400 ;
        RECT 487.5000 220.7550 489.5000 222.7550 ;
        RECT 479.3500 220.7550 481.3500 222.7550 ;
        RECT 471.2000 220.7550 473.2000 222.7550 ;
        RECT 463.0500 220.7550 465.0500 222.7550 ;
        RECT 487.5000 213.6600 489.5000 215.6600 ;
        RECT 479.3500 213.6600 481.3500 215.6600 ;
        RECT 471.2000 213.6600 473.2000 215.6600 ;
        RECT 463.0500 213.6600 465.0500 215.6600 ;
        RECT 471.2000 227.8500 473.2000 229.8500 ;
        RECT 463.0500 227.8500 465.0500 229.8500 ;
        RECT 479.3500 227.8500 481.3500 229.8500 ;
        RECT 487.5000 227.8500 489.5000 229.8500 ;
        RECT 463.0500 234.9450 465.0500 236.9450 ;
        RECT 471.2000 234.9450 473.2000 236.9450 ;
        RECT 479.3500 234.9450 481.3500 236.9450 ;
        RECT 487.5000 234.9450 489.5000 236.9450 ;
        RECT 463.0500 242.0400 465.0500 244.0400 ;
        RECT 471.2000 242.0400 473.2000 244.0400 ;
        RECT 479.3500 242.0400 481.3500 244.0400 ;
        RECT 487.5000 242.0400 489.5000 244.0400 ;
        RECT 454.9000 249.1350 456.9000 251.1350 ;
        RECT 454.9000 256.2300 456.9000 258.2300 ;
        RECT 454.9000 263.3250 456.9000 265.3250 ;
        RECT 454.9000 270.4200 456.9000 272.4200 ;
        RECT 454.9000 277.5150 456.9000 279.5150 ;
        RECT 446.7500 256.2300 448.7500 258.2300 ;
        RECT 438.6000 256.2300 440.6000 258.2300 ;
        RECT 430.4500 256.2300 432.4500 258.2300 ;
        RECT 422.3000 256.2300 424.3000 258.2300 ;
        RECT 446.7500 249.1350 448.7500 251.1350 ;
        RECT 438.6000 249.1350 440.6000 251.1350 ;
        RECT 430.4500 249.1350 432.4500 251.1350 ;
        RECT 422.3000 249.1350 424.3000 251.1350 ;
        RECT 430.4500 263.3250 432.4500 265.3250 ;
        RECT 422.3000 263.3250 424.3000 265.3250 ;
        RECT 438.6000 263.3250 440.6000 265.3250 ;
        RECT 446.7500 263.3250 448.7500 265.3250 ;
        RECT 422.3000 270.4200 424.3000 272.4200 ;
        RECT 430.4500 270.4200 432.4500 272.4200 ;
        RECT 438.6000 270.4200 440.6000 272.4200 ;
        RECT 446.7500 270.4200 448.7500 272.4200 ;
        RECT 422.3000 277.5150 424.3000 279.5150 ;
        RECT 430.4500 277.5150 432.4500 279.5150 ;
        RECT 438.6000 277.5150 440.6000 279.5150 ;
        RECT 446.7500 277.5150 448.7500 279.5150 ;
        RECT 487.5000 256.2300 489.5000 258.2300 ;
        RECT 479.3500 256.2300 481.3500 258.2300 ;
        RECT 471.2000 256.2300 473.2000 258.2300 ;
        RECT 463.0500 256.2300 465.0500 258.2300 ;
        RECT 487.5000 249.1350 489.5000 251.1350 ;
        RECT 479.3500 249.1350 481.3500 251.1350 ;
        RECT 471.2000 249.1350 473.2000 251.1350 ;
        RECT 463.0500 249.1350 465.0500 251.1350 ;
        RECT 471.2000 263.3250 473.2000 265.3250 ;
        RECT 463.0500 263.3250 465.0500 265.3250 ;
        RECT 479.3500 263.3250 481.3500 265.3250 ;
        RECT 487.5000 263.3250 489.5000 265.3250 ;
        RECT 463.0500 270.4200 465.0500 272.4200 ;
        RECT 471.2000 270.4200 473.2000 272.4200 ;
        RECT 479.3500 270.4200 481.3500 272.4200 ;
        RECT 487.5000 270.4200 489.5000 272.4200 ;
        RECT 463.0500 277.5150 465.0500 279.5150 ;
        RECT 471.2000 277.5150 473.2000 279.5150 ;
        RECT 479.3500 277.5150 481.3500 279.5150 ;
        RECT 487.5000 277.5150 489.5000 279.5150 ;
        RECT 520.1000 220.7550 522.1000 222.7550 ;
        RECT 511.9500 220.7550 513.9500 222.7550 ;
        RECT 503.8000 220.7550 505.8000 222.7550 ;
        RECT 495.6500 220.7550 497.6500 222.7550 ;
        RECT 520.1000 213.6600 522.1000 215.6600 ;
        RECT 511.9500 213.6600 513.9500 215.6600 ;
        RECT 503.8000 213.6600 505.8000 215.6600 ;
        RECT 495.6500 213.6600 497.6500 215.6600 ;
        RECT 503.8000 227.8500 505.8000 229.8500 ;
        RECT 495.6500 227.8500 497.6500 229.8500 ;
        RECT 511.9500 227.8500 513.9500 229.8500 ;
        RECT 520.1000 227.8500 522.1000 229.8500 ;
        RECT 495.6500 234.9450 497.6500 236.9450 ;
        RECT 503.8000 234.9450 505.8000 236.9450 ;
        RECT 511.9500 234.9450 513.9500 236.9450 ;
        RECT 520.1000 234.9450 522.1000 236.9450 ;
        RECT 495.6500 242.0400 497.6500 244.0400 ;
        RECT 503.8000 242.0400 505.8000 244.0400 ;
        RECT 511.9500 242.0400 513.9500 244.0400 ;
        RECT 520.1000 242.0400 522.1000 244.0400 ;
        RECT 552.7000 220.7550 554.7000 222.7550 ;
        RECT 544.5500 220.7550 546.5500 222.7550 ;
        RECT 536.4000 220.7550 538.4000 222.7550 ;
        RECT 528.2500 220.7550 530.2500 222.7550 ;
        RECT 552.7000 213.6600 554.7000 215.6600 ;
        RECT 544.5500 213.6600 546.5500 215.6600 ;
        RECT 536.4000 213.6600 538.4000 215.6600 ;
        RECT 528.2500 213.6600 530.2500 215.6600 ;
        RECT 536.4000 227.8500 538.4000 229.8500 ;
        RECT 528.2500 227.8500 530.2500 229.8500 ;
        RECT 544.5500 227.8500 546.5500 229.8500 ;
        RECT 552.7000 227.8500 554.7000 229.8500 ;
        RECT 528.2500 234.9450 530.2500 236.9450 ;
        RECT 536.4000 234.9450 538.4000 236.9450 ;
        RECT 544.5500 234.9450 546.5500 236.9450 ;
        RECT 552.7000 234.9450 554.7000 236.9450 ;
        RECT 528.2500 242.0400 530.2500 244.0400 ;
        RECT 536.4000 242.0400 538.4000 244.0400 ;
        RECT 544.5500 242.0400 546.5500 244.0400 ;
        RECT 552.7000 242.0400 554.7000 244.0400 ;
        RECT 520.1000 256.2300 522.1000 258.2300 ;
        RECT 511.9500 256.2300 513.9500 258.2300 ;
        RECT 503.8000 256.2300 505.8000 258.2300 ;
        RECT 495.6500 256.2300 497.6500 258.2300 ;
        RECT 520.1000 249.1350 522.1000 251.1350 ;
        RECT 511.9500 249.1350 513.9500 251.1350 ;
        RECT 503.8000 249.1350 505.8000 251.1350 ;
        RECT 495.6500 249.1350 497.6500 251.1350 ;
        RECT 503.8000 263.3250 505.8000 265.3250 ;
        RECT 495.6500 263.3250 497.6500 265.3250 ;
        RECT 511.9500 263.3250 513.9500 265.3250 ;
        RECT 520.1000 263.3250 522.1000 265.3250 ;
        RECT 495.6500 270.4200 497.6500 272.4200 ;
        RECT 503.8000 270.4200 505.8000 272.4200 ;
        RECT 511.9500 270.4200 513.9500 272.4200 ;
        RECT 520.1000 270.4200 522.1000 272.4200 ;
        RECT 495.6500 277.5150 497.6500 279.5150 ;
        RECT 503.8000 277.5150 505.8000 279.5150 ;
        RECT 511.9500 277.5150 513.9500 279.5150 ;
        RECT 520.1000 277.5150 522.1000 279.5150 ;
        RECT 552.7000 256.2300 554.7000 258.2300 ;
        RECT 544.5500 256.2300 546.5500 258.2300 ;
        RECT 536.4000 256.2300 538.4000 258.2300 ;
        RECT 528.2500 256.2300 530.2500 258.2300 ;
        RECT 552.7000 249.1350 554.7000 251.1350 ;
        RECT 544.5500 249.1350 546.5500 251.1350 ;
        RECT 536.4000 249.1350 538.4000 251.1350 ;
        RECT 528.2500 249.1350 530.2500 251.1350 ;
        RECT 536.4000 263.3250 538.4000 265.3250 ;
        RECT 528.2500 263.3250 530.2500 265.3250 ;
        RECT 544.5500 263.3250 546.5500 265.3250 ;
        RECT 552.7000 263.3250 554.7000 265.3250 ;
        RECT 528.2500 270.4200 530.2500 272.4200 ;
        RECT 536.4000 270.4200 538.4000 272.4200 ;
        RECT 544.5500 270.4200 546.5500 272.4200 ;
        RECT 552.7000 270.4200 554.7000 272.4200 ;
        RECT 528.2500 277.5150 530.2500 279.5150 ;
        RECT 536.4000 277.5150 538.4000 279.5150 ;
        RECT 544.5500 277.5150 546.5500 279.5150 ;
        RECT 552.7000 277.5150 554.7000 279.5150 ;
        RECT 6.0000 419.4150 8.0000 421.4150 ;
        RECT 44.0000 419.4150 46.0000 421.4150 ;
        RECT 60.0000 419.4150 62.0000 421.4150 ;
        RECT 68.5150 419.4150 70.5150 421.4150 ;
        RECT 77.0300 419.4150 79.0300 421.4150 ;
        RECT 85.5450 419.4150 87.5450 421.4150 ;
        RECT 94.0600 419.4150 96.0600 421.4150 ;
        RECT 102.5750 419.4150 104.5750 421.4150 ;
        RECT 111.0900 419.4150 113.0900 421.4150 ;
        RECT 119.6050 419.4150 121.6050 421.4150 ;
        RECT 128.1200 419.4150 130.1200 421.4150 ;
        RECT 136.6350 419.4150 138.6350 421.4150 ;
        RECT 204.7550 419.4150 206.7550 421.4150 ;
        RECT 196.2400 419.4150 198.2400 421.4150 ;
        RECT 187.7250 419.4150 189.7250 421.4150 ;
        RECT 179.2100 419.4150 181.2100 421.4150 ;
        RECT 170.6950 419.4150 172.6950 421.4150 ;
        RECT 162.1800 419.4150 164.1800 421.4150 ;
        RECT 153.6650 419.4150 155.6650 421.4150 ;
        RECT 145.1500 419.4150 147.1500 421.4150 ;
        RECT 255.8450 419.4150 257.8450 421.4150 ;
        RECT 247.3300 419.4150 249.3300 421.4150 ;
        RECT 238.8150 419.4150 240.8150 421.4150 ;
        RECT 230.3000 419.4150 232.3000 421.4150 ;
        RECT 221.7850 419.4150 223.7850 421.4150 ;
        RECT 213.2700 419.4150 215.2700 421.4150 ;
        RECT 264.3600 419.4150 266.3600 421.4150 ;
        RECT 272.8750 419.4150 274.8750 421.4150 ;
        RECT 6.0000 348.4650 8.0000 350.4650 ;
        RECT 68.5150 284.6100 70.5150 286.6100 ;
        RECT 68.5150 291.7050 70.5150 293.7050 ;
        RECT 68.5150 298.8000 70.5150 300.8000 ;
        RECT 68.5150 305.8950 70.5150 307.8950 ;
        RECT 68.5150 312.9900 70.5150 314.9900 ;
        RECT 68.5150 320.0850 70.5150 322.0850 ;
        RECT 68.5150 327.1800 70.5150 329.1800 ;
        RECT 6.0000 291.7050 8.0000 293.7050 ;
        RECT 6.0000 284.6100 8.0000 286.6100 ;
        RECT 6.0000 305.8950 8.0000 307.8950 ;
        RECT 6.0000 298.8000 8.0000 300.8000 ;
        RECT 6.0000 312.9900 8.0000 314.9900 ;
        RECT 44.0000 291.7050 46.0000 293.7050 ;
        RECT 44.0000 284.6100 46.0000 286.6100 ;
        RECT 60.0000 284.6100 62.0000 286.6100 ;
        RECT 60.0000 291.7050 62.0000 293.7050 ;
        RECT 44.0000 298.8000 46.0000 300.8000 ;
        RECT 44.0000 305.8950 46.0000 307.8950 ;
        RECT 44.0000 312.9900 46.0000 314.9900 ;
        RECT 60.0000 298.8000 62.0000 300.8000 ;
        RECT 60.0000 305.8950 62.0000 307.8950 ;
        RECT 60.0000 312.9900 62.0000 314.9900 ;
        RECT 6.0000 320.0850 8.0000 322.0850 ;
        RECT 6.0000 327.1800 8.0000 329.1800 ;
        RECT 6.0000 341.3700 8.0000 343.3700 ;
        RECT 6.0000 334.2750 8.0000 336.2750 ;
        RECT 44.0000 320.0850 46.0000 322.0850 ;
        RECT 44.0000 327.1800 46.0000 329.1800 ;
        RECT 60.0000 327.1800 62.0000 329.1800 ;
        RECT 60.0000 320.0850 62.0000 322.0850 ;
        RECT 44.0000 341.3700 46.0000 343.3700 ;
        RECT 44.0000 334.2750 46.0000 336.2750 ;
        RECT 102.5750 291.7050 104.5750 293.7050 ;
        RECT 94.0600 291.7050 96.0600 293.7050 ;
        RECT 85.5450 291.7050 87.5450 293.7050 ;
        RECT 77.0300 291.7050 79.0300 293.7050 ;
        RECT 102.5750 284.6100 104.5750 286.6100 ;
        RECT 94.0600 284.6100 96.0600 286.6100 ;
        RECT 85.5450 284.6100 87.5450 286.6100 ;
        RECT 77.0300 284.6100 79.0300 286.6100 ;
        RECT 85.5450 298.8000 87.5450 300.8000 ;
        RECT 77.0300 298.8000 79.0300 300.8000 ;
        RECT 94.0600 298.8000 96.0600 300.8000 ;
        RECT 102.5750 298.8000 104.5750 300.8000 ;
        RECT 77.0300 305.8950 79.0300 307.8950 ;
        RECT 85.5450 305.8950 87.5450 307.8950 ;
        RECT 94.0600 305.8950 96.0600 307.8950 ;
        RECT 102.5750 305.8950 104.5750 307.8950 ;
        RECT 77.0300 312.9900 79.0300 314.9900 ;
        RECT 85.5450 312.9900 87.5450 314.9900 ;
        RECT 94.0600 312.9900 96.0600 314.9900 ;
        RECT 102.5750 312.9900 104.5750 314.9900 ;
        RECT 136.6350 291.7050 138.6350 293.7050 ;
        RECT 128.1200 291.7050 130.1200 293.7050 ;
        RECT 119.6050 291.7050 121.6050 293.7050 ;
        RECT 111.0900 291.7050 113.0900 293.7050 ;
        RECT 136.6350 284.6100 138.6350 286.6100 ;
        RECT 128.1200 284.6100 130.1200 286.6100 ;
        RECT 119.6050 284.6100 121.6050 286.6100 ;
        RECT 111.0900 284.6100 113.0900 286.6100 ;
        RECT 119.6050 298.8000 121.6050 300.8000 ;
        RECT 111.0900 298.8000 113.0900 300.8000 ;
        RECT 128.1200 298.8000 130.1200 300.8000 ;
        RECT 136.6350 298.8000 138.6350 300.8000 ;
        RECT 111.0900 305.8950 113.0900 307.8950 ;
        RECT 119.6050 305.8950 121.6050 307.8950 ;
        RECT 128.1200 305.8950 130.1200 307.8950 ;
        RECT 136.6350 305.8950 138.6350 307.8950 ;
        RECT 111.0900 312.9900 113.0900 314.9900 ;
        RECT 119.6050 312.9900 121.6050 314.9900 ;
        RECT 128.1200 312.9900 130.1200 314.9900 ;
        RECT 136.6350 312.9900 138.6350 314.9900 ;
        RECT 102.5750 327.1800 104.5750 329.1800 ;
        RECT 94.0600 327.1800 96.0600 329.1800 ;
        RECT 85.5450 327.1800 87.5450 329.1800 ;
        RECT 77.0300 327.1800 79.0300 329.1800 ;
        RECT 102.5750 320.0850 104.5750 322.0850 ;
        RECT 94.0600 320.0850 96.0600 322.0850 ;
        RECT 85.5450 320.0850 87.5450 322.0850 ;
        RECT 77.0300 320.0850 79.0300 322.0850 ;
        RECT 119.6050 327.1800 121.6050 329.1800 ;
        RECT 111.0900 327.1800 113.0900 329.1800 ;
        RECT 136.6350 320.0850 138.6350 322.0850 ;
        RECT 128.1200 320.0850 130.1200 322.0850 ;
        RECT 119.6050 320.0850 121.6050 322.0850 ;
        RECT 111.0900 320.0850 113.0900 322.0850 ;
        RECT 128.1200 327.1800 130.1200 329.1800 ;
        RECT 136.6350 327.1800 138.6350 329.1800 ;
        RECT 68.5150 412.3200 70.5150 414.3200 ;
        RECT 6.0000 383.9400 8.0000 385.9400 ;
        RECT 6.0000 355.5600 8.0000 357.5600 ;
        RECT 6.0000 362.6550 8.0000 364.6550 ;
        RECT 6.0000 369.7500 8.0000 371.7500 ;
        RECT 6.0000 376.8450 8.0000 378.8450 ;
        RECT 6.0000 398.1300 8.0000 400.1300 ;
        RECT 6.0000 391.0350 8.0000 393.0350 ;
        RECT 6.0000 412.3200 8.0000 414.3200 ;
        RECT 6.0000 405.2250 8.0000 407.2250 ;
        RECT 44.0000 398.1300 46.0000 400.1300 ;
        RECT 44.0000 412.3200 46.0000 414.3200 ;
        RECT 44.0000 405.2250 46.0000 407.2250 ;
        RECT 60.0000 412.3200 62.0000 414.3200 ;
        RECT 77.0300 412.3200 79.0300 414.3200 ;
        RECT 85.5450 412.3200 87.5450 414.3200 ;
        RECT 94.0600 412.3200 96.0600 414.3200 ;
        RECT 102.5750 412.3200 104.5750 414.3200 ;
        RECT 111.0900 412.3200 113.0900 414.3200 ;
        RECT 119.6050 412.3200 121.6050 414.3200 ;
        RECT 128.1200 412.3200 130.1200 414.3200 ;
        RECT 136.6350 412.3200 138.6350 414.3200 ;
        RECT 170.6950 291.7050 172.6950 293.7050 ;
        RECT 162.1800 291.7050 164.1800 293.7050 ;
        RECT 153.6650 291.7050 155.6650 293.7050 ;
        RECT 145.1500 291.7050 147.1500 293.7050 ;
        RECT 170.6950 284.6100 172.6950 286.6100 ;
        RECT 162.1800 284.6100 164.1800 286.6100 ;
        RECT 153.6650 284.6100 155.6650 286.6100 ;
        RECT 145.1500 284.6100 147.1500 286.6100 ;
        RECT 153.6650 298.8000 155.6650 300.8000 ;
        RECT 145.1500 298.8000 147.1500 300.8000 ;
        RECT 162.1800 298.8000 164.1800 300.8000 ;
        RECT 170.6950 298.8000 172.6950 300.8000 ;
        RECT 145.1500 305.8950 147.1500 307.8950 ;
        RECT 153.6650 305.8950 155.6650 307.8950 ;
        RECT 162.1800 305.8950 164.1800 307.8950 ;
        RECT 170.6950 305.8950 172.6950 307.8950 ;
        RECT 145.1500 312.9900 147.1500 314.9900 ;
        RECT 153.6650 312.9900 155.6650 314.9900 ;
        RECT 162.1800 312.9900 164.1800 314.9900 ;
        RECT 170.6950 312.9900 172.6950 314.9900 ;
        RECT 204.7550 291.7050 206.7550 293.7050 ;
        RECT 196.2400 291.7050 198.2400 293.7050 ;
        RECT 187.7250 291.7050 189.7250 293.7050 ;
        RECT 179.2100 291.7050 181.2100 293.7050 ;
        RECT 204.7550 284.6100 206.7550 286.6100 ;
        RECT 196.2400 284.6100 198.2400 286.6100 ;
        RECT 187.7250 284.6100 189.7250 286.6100 ;
        RECT 179.2100 284.6100 181.2100 286.6100 ;
        RECT 187.7250 298.8000 189.7250 300.8000 ;
        RECT 179.2100 298.8000 181.2100 300.8000 ;
        RECT 196.2400 298.8000 198.2400 300.8000 ;
        RECT 204.7550 298.8000 206.7550 300.8000 ;
        RECT 179.2100 305.8950 181.2100 307.8950 ;
        RECT 187.7250 305.8950 189.7250 307.8950 ;
        RECT 196.2400 305.8950 198.2400 307.8950 ;
        RECT 204.7550 305.8950 206.7550 307.8950 ;
        RECT 179.2100 312.9900 181.2100 314.9900 ;
        RECT 187.7250 312.9900 189.7250 314.9900 ;
        RECT 196.2400 312.9900 198.2400 314.9900 ;
        RECT 204.7550 312.9900 206.7550 314.9900 ;
        RECT 170.6950 327.1800 172.6950 329.1800 ;
        RECT 162.1800 327.1800 164.1800 329.1800 ;
        RECT 153.6650 327.1800 155.6650 329.1800 ;
        RECT 145.1500 327.1800 147.1500 329.1800 ;
        RECT 170.6950 320.0850 172.6950 322.0850 ;
        RECT 162.1800 320.0850 164.1800 322.0850 ;
        RECT 153.6650 320.0850 155.6650 322.0850 ;
        RECT 145.1500 320.0850 147.1500 322.0850 ;
        RECT 187.7250 327.1800 189.7250 329.1800 ;
        RECT 179.2100 327.1800 181.2100 329.1800 ;
        RECT 204.7550 320.0850 206.7550 322.0850 ;
        RECT 196.2400 320.0850 198.2400 322.0850 ;
        RECT 187.7250 320.0850 189.7250 322.0850 ;
        RECT 179.2100 320.0850 181.2100 322.0850 ;
        RECT 196.2400 327.1800 198.2400 329.1800 ;
        RECT 204.7550 327.1800 206.7550 329.1800 ;
        RECT 238.8150 291.7050 240.8150 293.7050 ;
        RECT 230.3000 291.7050 232.3000 293.7050 ;
        RECT 221.7850 291.7050 223.7850 293.7050 ;
        RECT 213.2700 291.7050 215.2700 293.7050 ;
        RECT 238.8150 284.6100 240.8150 286.6100 ;
        RECT 230.3000 284.6100 232.3000 286.6100 ;
        RECT 221.7850 284.6100 223.7850 286.6100 ;
        RECT 213.2700 284.6100 215.2700 286.6100 ;
        RECT 221.7850 298.8000 223.7850 300.8000 ;
        RECT 213.2700 298.8000 215.2700 300.8000 ;
        RECT 230.3000 298.8000 232.3000 300.8000 ;
        RECT 238.8150 298.8000 240.8150 300.8000 ;
        RECT 213.2700 305.8950 215.2700 307.8950 ;
        RECT 221.7850 305.8950 223.7850 307.8950 ;
        RECT 230.3000 305.8950 232.3000 307.8950 ;
        RECT 238.8150 305.8950 240.8150 307.8950 ;
        RECT 213.2700 312.9900 215.2700 314.9900 ;
        RECT 221.7850 312.9900 223.7850 314.9900 ;
        RECT 230.3000 312.9900 232.3000 314.9900 ;
        RECT 238.8150 312.9900 240.8150 314.9900 ;
        RECT 272.8750 291.7050 274.8750 293.7050 ;
        RECT 264.3600 291.7050 266.3600 293.7050 ;
        RECT 255.8450 291.7050 257.8450 293.7050 ;
        RECT 247.3300 291.7050 249.3300 293.7050 ;
        RECT 272.8750 284.6100 274.8750 286.6100 ;
        RECT 264.3600 284.6100 266.3600 286.6100 ;
        RECT 255.8450 284.6100 257.8450 286.6100 ;
        RECT 247.3300 284.6100 249.3300 286.6100 ;
        RECT 255.8450 298.8000 257.8450 300.8000 ;
        RECT 247.3300 298.8000 249.3300 300.8000 ;
        RECT 264.3600 298.8000 266.3600 300.8000 ;
        RECT 272.8750 298.8000 274.8750 300.8000 ;
        RECT 247.3300 305.8950 249.3300 307.8950 ;
        RECT 255.8450 305.8950 257.8450 307.8950 ;
        RECT 264.3600 305.8950 266.3600 307.8950 ;
        RECT 272.8750 305.8950 274.8750 307.8950 ;
        RECT 247.3300 312.9900 249.3300 314.9900 ;
        RECT 255.8450 312.9900 257.8450 314.9900 ;
        RECT 264.3600 312.9900 266.3600 314.9900 ;
        RECT 272.8750 312.9900 274.8750 314.9900 ;
        RECT 238.8150 327.1800 240.8150 329.1800 ;
        RECT 230.3000 327.1800 232.3000 329.1800 ;
        RECT 221.7850 327.1800 223.7850 329.1800 ;
        RECT 213.2700 327.1800 215.2700 329.1800 ;
        RECT 238.8150 320.0850 240.8150 322.0850 ;
        RECT 230.3000 320.0850 232.3000 322.0850 ;
        RECT 221.7850 320.0850 223.7850 322.0850 ;
        RECT 213.2700 320.0850 215.2700 322.0850 ;
        RECT 255.8450 327.1800 257.8450 329.1800 ;
        RECT 247.3300 327.1800 249.3300 329.1800 ;
        RECT 272.8750 320.0850 274.8750 322.0850 ;
        RECT 264.3600 320.0850 266.3600 322.0850 ;
        RECT 255.8450 320.0850 257.8450 322.0850 ;
        RECT 247.3300 320.0850 249.3300 322.0850 ;
        RECT 264.3600 327.1800 266.3600 329.1800 ;
        RECT 272.8750 327.1800 274.8750 329.1800 ;
        RECT 204.7550 412.3200 206.7550 414.3200 ;
        RECT 196.2400 412.3200 198.2400 414.3200 ;
        RECT 187.7250 412.3200 189.7250 414.3200 ;
        RECT 179.2100 412.3200 181.2100 414.3200 ;
        RECT 170.6950 412.3200 172.6950 414.3200 ;
        RECT 162.1800 412.3200 164.1800 414.3200 ;
        RECT 153.6650 412.3200 155.6650 414.3200 ;
        RECT 145.1500 412.3200 147.1500 414.3200 ;
        RECT 255.8450 412.3200 257.8450 414.3200 ;
        RECT 247.3300 412.3200 249.3300 414.3200 ;
        RECT 238.8150 412.3200 240.8150 414.3200 ;
        RECT 230.3000 412.3200 232.3000 414.3200 ;
        RECT 221.7850 412.3200 223.7850 414.3200 ;
        RECT 213.2700 412.3200 215.2700 414.3200 ;
        RECT 264.3600 412.3200 266.3600 414.3200 ;
        RECT 272.8750 412.3200 274.8750 414.3200 ;
        RECT 68.5150 426.5100 70.5150 428.5100 ;
        RECT 68.5150 433.6050 70.5150 435.6050 ;
        RECT 68.5150 440.7000 70.5150 442.7000 ;
        RECT 68.5150 447.7950 70.5150 449.7950 ;
        RECT 68.5150 454.8900 70.5150 456.8900 ;
        RECT 68.5150 461.9850 70.5150 463.9850 ;
        RECT 68.5150 469.0800 70.5150 471.0800 ;
        RECT 68.5150 476.1750 70.5150 478.1750 ;
        RECT 68.5150 483.2700 70.5150 485.2700 ;
        RECT 44.0000 454.8900 46.0000 456.8900 ;
        RECT 6.0000 454.8900 8.0000 456.8900 ;
        RECT 60.0000 454.8900 62.0000 456.8900 ;
        RECT 6.0000 426.5100 8.0000 428.5100 ;
        RECT 6.0000 433.6050 8.0000 435.6050 ;
        RECT 6.0000 440.7000 8.0000 442.7000 ;
        RECT 6.0000 447.7950 8.0000 449.7950 ;
        RECT 44.0000 426.5100 46.0000 428.5100 ;
        RECT 44.0000 433.6050 46.0000 435.6050 ;
        RECT 60.0000 433.6050 62.0000 435.6050 ;
        RECT 60.0000 426.5100 62.0000 428.5100 ;
        RECT 44.0000 440.7000 46.0000 442.7000 ;
        RECT 44.0000 447.7950 46.0000 449.7950 ;
        RECT 60.0000 447.7950 62.0000 449.7950 ;
        RECT 60.0000 440.7000 62.0000 442.7000 ;
        RECT 6.0000 469.0800 8.0000 471.0800 ;
        RECT 6.0000 461.9850 8.0000 463.9850 ;
        RECT 6.0000 483.2700 8.0000 485.2700 ;
        RECT 6.0000 476.1750 8.0000 478.1750 ;
        RECT 44.0000 469.0800 46.0000 471.0800 ;
        RECT 44.0000 461.9850 46.0000 463.9850 ;
        RECT 60.0000 461.9850 62.0000 463.9850 ;
        RECT 60.0000 469.0800 62.0000 471.0800 ;
        RECT 44.0000 483.2700 46.0000 485.2700 ;
        RECT 44.0000 476.1750 46.0000 478.1750 ;
        RECT 60.0000 476.1750 62.0000 478.1750 ;
        RECT 60.0000 483.2700 62.0000 485.2700 ;
        RECT 77.0300 454.8900 79.0300 456.8900 ;
        RECT 85.5450 454.8900 87.5450 456.8900 ;
        RECT 94.0600 454.8900 96.0600 456.8900 ;
        RECT 102.5750 454.8900 104.5750 456.8900 ;
        RECT 111.0900 454.8900 113.0900 456.8900 ;
        RECT 119.6050 454.8900 121.6050 456.8900 ;
        RECT 128.1200 454.8900 130.1200 456.8900 ;
        RECT 136.6350 454.8900 138.6350 456.8900 ;
        RECT 102.5750 433.6050 104.5750 435.6050 ;
        RECT 94.0600 433.6050 96.0600 435.6050 ;
        RECT 85.5450 433.6050 87.5450 435.6050 ;
        RECT 77.0300 433.6050 79.0300 435.6050 ;
        RECT 102.5750 426.5100 104.5750 428.5100 ;
        RECT 94.0600 426.5100 96.0600 428.5100 ;
        RECT 85.5450 426.5100 87.5450 428.5100 ;
        RECT 77.0300 426.5100 79.0300 428.5100 ;
        RECT 85.5450 447.7950 87.5450 449.7950 ;
        RECT 77.0300 447.7950 79.0300 449.7950 ;
        RECT 102.5750 440.7000 104.5750 442.7000 ;
        RECT 94.0600 440.7000 96.0600 442.7000 ;
        RECT 85.5450 440.7000 87.5450 442.7000 ;
        RECT 77.0300 440.7000 79.0300 442.7000 ;
        RECT 94.0600 447.7950 96.0600 449.7950 ;
        RECT 102.5750 447.7950 104.5750 449.7950 ;
        RECT 136.6350 433.6050 138.6350 435.6050 ;
        RECT 128.1200 433.6050 130.1200 435.6050 ;
        RECT 119.6050 433.6050 121.6050 435.6050 ;
        RECT 111.0900 433.6050 113.0900 435.6050 ;
        RECT 136.6350 426.5100 138.6350 428.5100 ;
        RECT 128.1200 426.5100 130.1200 428.5100 ;
        RECT 119.6050 426.5100 121.6050 428.5100 ;
        RECT 111.0900 426.5100 113.0900 428.5100 ;
        RECT 119.6050 447.7950 121.6050 449.7950 ;
        RECT 111.0900 447.7950 113.0900 449.7950 ;
        RECT 136.6350 440.7000 138.6350 442.7000 ;
        RECT 128.1200 440.7000 130.1200 442.7000 ;
        RECT 119.6050 440.7000 121.6050 442.7000 ;
        RECT 111.0900 440.7000 113.0900 442.7000 ;
        RECT 128.1200 447.7950 130.1200 449.7950 ;
        RECT 136.6350 447.7950 138.6350 449.7950 ;
        RECT 102.5750 469.0800 104.5750 471.0800 ;
        RECT 94.0600 469.0800 96.0600 471.0800 ;
        RECT 85.5450 469.0800 87.5450 471.0800 ;
        RECT 77.0300 469.0800 79.0300 471.0800 ;
        RECT 102.5750 461.9850 104.5750 463.9850 ;
        RECT 94.0600 461.9850 96.0600 463.9850 ;
        RECT 85.5450 461.9850 87.5450 463.9850 ;
        RECT 77.0300 461.9850 79.0300 463.9850 ;
        RECT 85.5450 483.2700 87.5450 485.2700 ;
        RECT 77.0300 483.2700 79.0300 485.2700 ;
        RECT 102.5750 476.1750 104.5750 478.1750 ;
        RECT 94.0600 476.1750 96.0600 478.1750 ;
        RECT 85.5450 476.1750 87.5450 478.1750 ;
        RECT 77.0300 476.1750 79.0300 478.1750 ;
        RECT 94.0600 483.2700 96.0600 485.2700 ;
        RECT 102.5750 483.2700 104.5750 485.2700 ;
        RECT 136.6350 469.0800 138.6350 471.0800 ;
        RECT 128.1200 469.0800 130.1200 471.0800 ;
        RECT 119.6050 469.0800 121.6050 471.0800 ;
        RECT 111.0900 469.0800 113.0900 471.0800 ;
        RECT 136.6350 461.9850 138.6350 463.9850 ;
        RECT 128.1200 461.9850 130.1200 463.9850 ;
        RECT 119.6050 461.9850 121.6050 463.9850 ;
        RECT 111.0900 461.9850 113.0900 463.9850 ;
        RECT 119.6050 483.2700 121.6050 485.2700 ;
        RECT 111.0900 483.2700 113.0900 485.2700 ;
        RECT 136.6350 476.1750 138.6350 478.1750 ;
        RECT 128.1200 476.1750 130.1200 478.1750 ;
        RECT 119.6050 476.1750 121.6050 478.1750 ;
        RECT 111.0900 476.1750 113.0900 478.1750 ;
        RECT 128.1200 483.2700 130.1200 485.2700 ;
        RECT 136.6350 483.2700 138.6350 485.2700 ;
        RECT 68.5150 490.3650 70.5150 492.3650 ;
        RECT 68.5150 497.4600 70.5150 499.4600 ;
        RECT 68.5150 504.5550 70.5150 506.5550 ;
        RECT 68.5150 511.6500 70.5150 513.6500 ;
        RECT 68.5150 518.7450 70.5150 520.7450 ;
        RECT 68.5150 525.8400 70.5150 527.8400 ;
        RECT 68.5150 532.9350 70.5150 534.9350 ;
        RECT 68.5150 540.0300 70.5150 542.0300 ;
        RECT 68.5150 547.1250 70.5150 549.1250 ;
        RECT 68.5150 554.2200 70.5150 556.2200 ;
        RECT 6.0000 497.4600 8.0000 499.4600 ;
        RECT 6.0000 490.3650 8.0000 492.3650 ;
        RECT 6.0000 504.5550 8.0000 506.5550 ;
        RECT 6.0000 511.6500 8.0000 513.6500 ;
        RECT 6.0000 518.7450 8.0000 520.7450 ;
        RECT 44.0000 490.3650 46.0000 492.3650 ;
        RECT 44.0000 497.4600 46.0000 499.4600 ;
        RECT 44.0000 504.5550 46.0000 506.5550 ;
        RECT 60.0000 490.3650 62.0000 492.3650 ;
        RECT 60.0000 497.4600 62.0000 499.4600 ;
        RECT 60.0000 504.5550 62.0000 506.5550 ;
        RECT 44.0000 511.6500 46.0000 513.6500 ;
        RECT 44.0000 518.7450 46.0000 520.7450 ;
        RECT 60.0000 518.7450 62.0000 520.7450 ;
        RECT 60.0000 511.6500 62.0000 513.6500 ;
        RECT 6.0000 532.9350 8.0000 534.9350 ;
        RECT 6.0000 525.8400 8.0000 527.8400 ;
        RECT 6.0000 540.0300 8.0000 542.0300 ;
        RECT 6.0000 547.1250 8.0000 549.1250 ;
        RECT 6.0000 554.2200 8.0000 556.2200 ;
        RECT 44.0000 525.8400 46.0000 527.8400 ;
        RECT 44.0000 532.9350 46.0000 534.9350 ;
        RECT 44.0000 540.0300 46.0000 542.0300 ;
        RECT 60.0000 532.9350 62.0000 534.9350 ;
        RECT 60.0000 525.8400 62.0000 527.8400 ;
        RECT 60.0000 540.0300 62.0000 542.0300 ;
        RECT 44.0000 547.1250 46.0000 549.1250 ;
        RECT 44.0000 554.2200 46.0000 556.2200 ;
        RECT 60.0000 554.2200 62.0000 556.2200 ;
        RECT 60.0000 547.1250 62.0000 549.1250 ;
        RECT 85.5450 504.5550 87.5450 506.5550 ;
        RECT 77.0300 504.5550 79.0300 506.5550 ;
        RECT 102.5750 497.4600 104.5750 499.4600 ;
        RECT 94.0600 497.4600 96.0600 499.4600 ;
        RECT 85.5450 497.4600 87.5450 499.4600 ;
        RECT 77.0300 497.4600 79.0300 499.4600 ;
        RECT 102.5750 490.3650 104.5750 492.3650 ;
        RECT 94.0600 490.3650 96.0600 492.3650 ;
        RECT 85.5450 490.3650 87.5450 492.3650 ;
        RECT 77.0300 490.3650 79.0300 492.3650 ;
        RECT 94.0600 504.5550 96.0600 506.5550 ;
        RECT 102.5750 504.5550 104.5750 506.5550 ;
        RECT 77.0300 511.6500 79.0300 513.6500 ;
        RECT 85.5450 511.6500 87.5450 513.6500 ;
        RECT 94.0600 511.6500 96.0600 513.6500 ;
        RECT 102.5750 511.6500 104.5750 513.6500 ;
        RECT 77.0300 518.7450 79.0300 520.7450 ;
        RECT 85.5450 518.7450 87.5450 520.7450 ;
        RECT 94.0600 518.7450 96.0600 520.7450 ;
        RECT 102.5750 518.7450 104.5750 520.7450 ;
        RECT 119.6050 504.5550 121.6050 506.5550 ;
        RECT 111.0900 504.5550 113.0900 506.5550 ;
        RECT 136.6350 497.4600 138.6350 499.4600 ;
        RECT 128.1200 497.4600 130.1200 499.4600 ;
        RECT 119.6050 497.4600 121.6050 499.4600 ;
        RECT 111.0900 497.4600 113.0900 499.4600 ;
        RECT 136.6350 490.3650 138.6350 492.3650 ;
        RECT 128.1200 490.3650 130.1200 492.3650 ;
        RECT 119.6050 490.3650 121.6050 492.3650 ;
        RECT 111.0900 490.3650 113.0900 492.3650 ;
        RECT 128.1200 504.5550 130.1200 506.5550 ;
        RECT 136.6350 504.5550 138.6350 506.5550 ;
        RECT 111.0900 511.6500 113.0900 513.6500 ;
        RECT 119.6050 511.6500 121.6050 513.6500 ;
        RECT 128.1200 511.6500 130.1200 513.6500 ;
        RECT 136.6350 511.6500 138.6350 513.6500 ;
        RECT 111.0900 518.7450 113.0900 520.7450 ;
        RECT 119.6050 518.7450 121.6050 520.7450 ;
        RECT 128.1200 518.7450 130.1200 520.7450 ;
        RECT 136.6350 518.7450 138.6350 520.7450 ;
        RECT 85.5450 540.0300 87.5450 542.0300 ;
        RECT 77.0300 540.0300 79.0300 542.0300 ;
        RECT 102.5750 532.9350 104.5750 534.9350 ;
        RECT 94.0600 532.9350 96.0600 534.9350 ;
        RECT 85.5450 532.9350 87.5450 534.9350 ;
        RECT 77.0300 532.9350 79.0300 534.9350 ;
        RECT 102.5750 525.8400 104.5750 527.8400 ;
        RECT 94.0600 525.8400 96.0600 527.8400 ;
        RECT 85.5450 525.8400 87.5450 527.8400 ;
        RECT 77.0300 525.8400 79.0300 527.8400 ;
        RECT 94.0600 540.0300 96.0600 542.0300 ;
        RECT 102.5750 540.0300 104.5750 542.0300 ;
        RECT 77.0300 547.1250 79.0300 549.1250 ;
        RECT 85.5450 547.1250 87.5450 549.1250 ;
        RECT 94.0600 547.1250 96.0600 549.1250 ;
        RECT 102.5750 547.1250 104.5750 549.1250 ;
        RECT 77.0300 554.2200 79.0300 556.2200 ;
        RECT 85.5450 554.2200 87.5450 556.2200 ;
        RECT 94.0600 554.2200 96.0600 556.2200 ;
        RECT 102.5750 554.2200 104.5750 556.2200 ;
        RECT 119.6050 540.0300 121.6050 542.0300 ;
        RECT 111.0900 540.0300 113.0900 542.0300 ;
        RECT 136.6350 532.9350 138.6350 534.9350 ;
        RECT 128.1200 532.9350 130.1200 534.9350 ;
        RECT 119.6050 532.9350 121.6050 534.9350 ;
        RECT 111.0900 532.9350 113.0900 534.9350 ;
        RECT 136.6350 525.8400 138.6350 527.8400 ;
        RECT 128.1200 525.8400 130.1200 527.8400 ;
        RECT 119.6050 525.8400 121.6050 527.8400 ;
        RECT 111.0900 525.8400 113.0900 527.8400 ;
        RECT 128.1200 540.0300 130.1200 542.0300 ;
        RECT 136.6350 540.0300 138.6350 542.0300 ;
        RECT 111.0900 547.1250 113.0900 549.1250 ;
        RECT 119.6050 547.1250 121.6050 549.1250 ;
        RECT 128.1200 547.1250 130.1200 549.1250 ;
        RECT 136.6350 547.1250 138.6350 549.1250 ;
        RECT 111.0900 554.2200 113.0900 556.2200 ;
        RECT 119.6050 554.2200 121.6050 556.2200 ;
        RECT 128.1200 554.2200 130.1200 556.2200 ;
        RECT 136.6350 554.2200 138.6350 556.2200 ;
        RECT 145.1500 454.8900 147.1500 456.8900 ;
        RECT 153.6650 454.8900 155.6650 456.8900 ;
        RECT 162.1800 454.8900 164.1800 456.8900 ;
        RECT 170.6950 454.8900 172.6950 456.8900 ;
        RECT 179.2100 454.8900 181.2100 456.8900 ;
        RECT 187.7250 454.8900 189.7250 456.8900 ;
        RECT 196.2400 454.8900 198.2400 456.8900 ;
        RECT 204.7550 454.8900 206.7550 456.8900 ;
        RECT 170.6950 433.6050 172.6950 435.6050 ;
        RECT 162.1800 433.6050 164.1800 435.6050 ;
        RECT 153.6650 433.6050 155.6650 435.6050 ;
        RECT 145.1500 433.6050 147.1500 435.6050 ;
        RECT 170.6950 426.5100 172.6950 428.5100 ;
        RECT 162.1800 426.5100 164.1800 428.5100 ;
        RECT 153.6650 426.5100 155.6650 428.5100 ;
        RECT 145.1500 426.5100 147.1500 428.5100 ;
        RECT 153.6650 447.7950 155.6650 449.7950 ;
        RECT 145.1500 447.7950 147.1500 449.7950 ;
        RECT 170.6950 440.7000 172.6950 442.7000 ;
        RECT 162.1800 440.7000 164.1800 442.7000 ;
        RECT 153.6650 440.7000 155.6650 442.7000 ;
        RECT 145.1500 440.7000 147.1500 442.7000 ;
        RECT 162.1800 447.7950 164.1800 449.7950 ;
        RECT 170.6950 447.7950 172.6950 449.7950 ;
        RECT 204.7550 433.6050 206.7550 435.6050 ;
        RECT 196.2400 433.6050 198.2400 435.6050 ;
        RECT 187.7250 433.6050 189.7250 435.6050 ;
        RECT 179.2100 433.6050 181.2100 435.6050 ;
        RECT 204.7550 426.5100 206.7550 428.5100 ;
        RECT 196.2400 426.5100 198.2400 428.5100 ;
        RECT 187.7250 426.5100 189.7250 428.5100 ;
        RECT 179.2100 426.5100 181.2100 428.5100 ;
        RECT 187.7250 447.7950 189.7250 449.7950 ;
        RECT 179.2100 447.7950 181.2100 449.7950 ;
        RECT 204.7550 440.7000 206.7550 442.7000 ;
        RECT 196.2400 440.7000 198.2400 442.7000 ;
        RECT 187.7250 440.7000 189.7250 442.7000 ;
        RECT 179.2100 440.7000 181.2100 442.7000 ;
        RECT 196.2400 447.7950 198.2400 449.7950 ;
        RECT 204.7550 447.7950 206.7550 449.7950 ;
        RECT 170.6950 469.0800 172.6950 471.0800 ;
        RECT 162.1800 469.0800 164.1800 471.0800 ;
        RECT 153.6650 469.0800 155.6650 471.0800 ;
        RECT 145.1500 469.0800 147.1500 471.0800 ;
        RECT 170.6950 461.9850 172.6950 463.9850 ;
        RECT 162.1800 461.9850 164.1800 463.9850 ;
        RECT 153.6650 461.9850 155.6650 463.9850 ;
        RECT 145.1500 461.9850 147.1500 463.9850 ;
        RECT 153.6650 483.2700 155.6650 485.2700 ;
        RECT 145.1500 483.2700 147.1500 485.2700 ;
        RECT 170.6950 476.1750 172.6950 478.1750 ;
        RECT 162.1800 476.1750 164.1800 478.1750 ;
        RECT 153.6650 476.1750 155.6650 478.1750 ;
        RECT 145.1500 476.1750 147.1500 478.1750 ;
        RECT 162.1800 483.2700 164.1800 485.2700 ;
        RECT 170.6950 483.2700 172.6950 485.2700 ;
        RECT 204.7550 469.0800 206.7550 471.0800 ;
        RECT 196.2400 469.0800 198.2400 471.0800 ;
        RECT 187.7250 469.0800 189.7250 471.0800 ;
        RECT 179.2100 469.0800 181.2100 471.0800 ;
        RECT 204.7550 461.9850 206.7550 463.9850 ;
        RECT 196.2400 461.9850 198.2400 463.9850 ;
        RECT 187.7250 461.9850 189.7250 463.9850 ;
        RECT 179.2100 461.9850 181.2100 463.9850 ;
        RECT 187.7250 483.2700 189.7250 485.2700 ;
        RECT 179.2100 483.2700 181.2100 485.2700 ;
        RECT 204.7550 476.1750 206.7550 478.1750 ;
        RECT 196.2400 476.1750 198.2400 478.1750 ;
        RECT 187.7250 476.1750 189.7250 478.1750 ;
        RECT 179.2100 476.1750 181.2100 478.1750 ;
        RECT 196.2400 483.2700 198.2400 485.2700 ;
        RECT 204.7550 483.2700 206.7550 485.2700 ;
        RECT 213.2700 454.8900 215.2700 456.8900 ;
        RECT 221.7850 454.8900 223.7850 456.8900 ;
        RECT 230.3000 454.8900 232.3000 456.8900 ;
        RECT 238.8150 454.8900 240.8150 456.8900 ;
        RECT 247.3300 454.8900 249.3300 456.8900 ;
        RECT 255.8450 454.8900 257.8450 456.8900 ;
        RECT 264.3600 454.8900 266.3600 456.8900 ;
        RECT 272.8750 454.8900 274.8750 456.8900 ;
        RECT 238.8150 433.6050 240.8150 435.6050 ;
        RECT 230.3000 433.6050 232.3000 435.6050 ;
        RECT 221.7850 433.6050 223.7850 435.6050 ;
        RECT 213.2700 433.6050 215.2700 435.6050 ;
        RECT 238.8150 426.5100 240.8150 428.5100 ;
        RECT 230.3000 426.5100 232.3000 428.5100 ;
        RECT 221.7850 426.5100 223.7850 428.5100 ;
        RECT 213.2700 426.5100 215.2700 428.5100 ;
        RECT 221.7850 447.7950 223.7850 449.7950 ;
        RECT 213.2700 447.7950 215.2700 449.7950 ;
        RECT 238.8150 440.7000 240.8150 442.7000 ;
        RECT 230.3000 440.7000 232.3000 442.7000 ;
        RECT 221.7850 440.7000 223.7850 442.7000 ;
        RECT 213.2700 440.7000 215.2700 442.7000 ;
        RECT 230.3000 447.7950 232.3000 449.7950 ;
        RECT 238.8150 447.7950 240.8150 449.7950 ;
        RECT 272.8750 433.6050 274.8750 435.6050 ;
        RECT 264.3600 433.6050 266.3600 435.6050 ;
        RECT 255.8450 433.6050 257.8450 435.6050 ;
        RECT 247.3300 433.6050 249.3300 435.6050 ;
        RECT 272.8750 426.5100 274.8750 428.5100 ;
        RECT 264.3600 426.5100 266.3600 428.5100 ;
        RECT 255.8450 426.5100 257.8450 428.5100 ;
        RECT 247.3300 426.5100 249.3300 428.5100 ;
        RECT 255.8450 447.7950 257.8450 449.7950 ;
        RECT 247.3300 447.7950 249.3300 449.7950 ;
        RECT 272.8750 440.7000 274.8750 442.7000 ;
        RECT 264.3600 440.7000 266.3600 442.7000 ;
        RECT 255.8450 440.7000 257.8450 442.7000 ;
        RECT 247.3300 440.7000 249.3300 442.7000 ;
        RECT 264.3600 447.7950 266.3600 449.7950 ;
        RECT 272.8750 447.7950 274.8750 449.7950 ;
        RECT 238.8150 469.0800 240.8150 471.0800 ;
        RECT 230.3000 469.0800 232.3000 471.0800 ;
        RECT 221.7850 469.0800 223.7850 471.0800 ;
        RECT 213.2700 469.0800 215.2700 471.0800 ;
        RECT 238.8150 461.9850 240.8150 463.9850 ;
        RECT 230.3000 461.9850 232.3000 463.9850 ;
        RECT 221.7850 461.9850 223.7850 463.9850 ;
        RECT 213.2700 461.9850 215.2700 463.9850 ;
        RECT 221.7850 483.2700 223.7850 485.2700 ;
        RECT 213.2700 483.2700 215.2700 485.2700 ;
        RECT 238.8150 476.1750 240.8150 478.1750 ;
        RECT 230.3000 476.1750 232.3000 478.1750 ;
        RECT 221.7850 476.1750 223.7850 478.1750 ;
        RECT 213.2700 476.1750 215.2700 478.1750 ;
        RECT 230.3000 483.2700 232.3000 485.2700 ;
        RECT 238.8150 483.2700 240.8150 485.2700 ;
        RECT 272.8750 469.0800 274.8750 471.0800 ;
        RECT 264.3600 469.0800 266.3600 471.0800 ;
        RECT 255.8450 469.0800 257.8450 471.0800 ;
        RECT 247.3300 469.0800 249.3300 471.0800 ;
        RECT 272.8750 461.9850 274.8750 463.9850 ;
        RECT 264.3600 461.9850 266.3600 463.9850 ;
        RECT 255.8450 461.9850 257.8450 463.9850 ;
        RECT 247.3300 461.9850 249.3300 463.9850 ;
        RECT 255.8450 483.2700 257.8450 485.2700 ;
        RECT 247.3300 483.2700 249.3300 485.2700 ;
        RECT 272.8750 476.1750 274.8750 478.1750 ;
        RECT 264.3600 476.1750 266.3600 478.1750 ;
        RECT 255.8450 476.1750 257.8450 478.1750 ;
        RECT 247.3300 476.1750 249.3300 478.1750 ;
        RECT 264.3600 483.2700 266.3600 485.2700 ;
        RECT 272.8750 483.2700 274.8750 485.2700 ;
        RECT 153.6650 504.5550 155.6650 506.5550 ;
        RECT 145.1500 504.5550 147.1500 506.5550 ;
        RECT 170.6950 497.4600 172.6950 499.4600 ;
        RECT 162.1800 497.4600 164.1800 499.4600 ;
        RECT 153.6650 497.4600 155.6650 499.4600 ;
        RECT 145.1500 497.4600 147.1500 499.4600 ;
        RECT 170.6950 490.3650 172.6950 492.3650 ;
        RECT 162.1800 490.3650 164.1800 492.3650 ;
        RECT 153.6650 490.3650 155.6650 492.3650 ;
        RECT 145.1500 490.3650 147.1500 492.3650 ;
        RECT 162.1800 504.5550 164.1800 506.5550 ;
        RECT 170.6950 504.5550 172.6950 506.5550 ;
        RECT 145.1500 511.6500 147.1500 513.6500 ;
        RECT 153.6650 511.6500 155.6650 513.6500 ;
        RECT 162.1800 511.6500 164.1800 513.6500 ;
        RECT 170.6950 511.6500 172.6950 513.6500 ;
        RECT 145.1500 518.7450 147.1500 520.7450 ;
        RECT 153.6650 518.7450 155.6650 520.7450 ;
        RECT 162.1800 518.7450 164.1800 520.7450 ;
        RECT 170.6950 518.7450 172.6950 520.7450 ;
        RECT 187.7250 504.5550 189.7250 506.5550 ;
        RECT 179.2100 504.5550 181.2100 506.5550 ;
        RECT 204.7550 497.4600 206.7550 499.4600 ;
        RECT 196.2400 497.4600 198.2400 499.4600 ;
        RECT 187.7250 497.4600 189.7250 499.4600 ;
        RECT 179.2100 497.4600 181.2100 499.4600 ;
        RECT 204.7550 490.3650 206.7550 492.3650 ;
        RECT 196.2400 490.3650 198.2400 492.3650 ;
        RECT 187.7250 490.3650 189.7250 492.3650 ;
        RECT 179.2100 490.3650 181.2100 492.3650 ;
        RECT 196.2400 504.5550 198.2400 506.5550 ;
        RECT 204.7550 504.5550 206.7550 506.5550 ;
        RECT 179.2100 511.6500 181.2100 513.6500 ;
        RECT 187.7250 511.6500 189.7250 513.6500 ;
        RECT 196.2400 511.6500 198.2400 513.6500 ;
        RECT 204.7550 511.6500 206.7550 513.6500 ;
        RECT 179.2100 518.7450 181.2100 520.7450 ;
        RECT 187.7250 518.7450 189.7250 520.7450 ;
        RECT 196.2400 518.7450 198.2400 520.7450 ;
        RECT 204.7550 518.7450 206.7550 520.7450 ;
        RECT 153.6650 540.0300 155.6650 542.0300 ;
        RECT 145.1500 540.0300 147.1500 542.0300 ;
        RECT 170.6950 532.9350 172.6950 534.9350 ;
        RECT 162.1800 532.9350 164.1800 534.9350 ;
        RECT 153.6650 532.9350 155.6650 534.9350 ;
        RECT 145.1500 532.9350 147.1500 534.9350 ;
        RECT 170.6950 525.8400 172.6950 527.8400 ;
        RECT 162.1800 525.8400 164.1800 527.8400 ;
        RECT 153.6650 525.8400 155.6650 527.8400 ;
        RECT 145.1500 525.8400 147.1500 527.8400 ;
        RECT 162.1800 540.0300 164.1800 542.0300 ;
        RECT 170.6950 540.0300 172.6950 542.0300 ;
        RECT 145.1500 547.1250 147.1500 549.1250 ;
        RECT 153.6650 547.1250 155.6650 549.1250 ;
        RECT 162.1800 547.1250 164.1800 549.1250 ;
        RECT 170.6950 547.1250 172.6950 549.1250 ;
        RECT 145.1500 554.2200 147.1500 556.2200 ;
        RECT 153.6650 554.2200 155.6650 556.2200 ;
        RECT 162.1800 554.2200 164.1800 556.2200 ;
        RECT 170.6950 554.2200 172.6950 556.2200 ;
        RECT 187.7250 540.0300 189.7250 542.0300 ;
        RECT 179.2100 540.0300 181.2100 542.0300 ;
        RECT 204.7550 532.9350 206.7550 534.9350 ;
        RECT 196.2400 532.9350 198.2400 534.9350 ;
        RECT 187.7250 532.9350 189.7250 534.9350 ;
        RECT 179.2100 532.9350 181.2100 534.9350 ;
        RECT 204.7550 525.8400 206.7550 527.8400 ;
        RECT 196.2400 525.8400 198.2400 527.8400 ;
        RECT 187.7250 525.8400 189.7250 527.8400 ;
        RECT 179.2100 525.8400 181.2100 527.8400 ;
        RECT 196.2400 540.0300 198.2400 542.0300 ;
        RECT 204.7550 540.0300 206.7550 542.0300 ;
        RECT 179.2100 547.1250 181.2100 549.1250 ;
        RECT 187.7250 547.1250 189.7250 549.1250 ;
        RECT 196.2400 547.1250 198.2400 549.1250 ;
        RECT 204.7550 547.1250 206.7550 549.1250 ;
        RECT 179.2100 554.2200 181.2100 556.2200 ;
        RECT 187.7250 554.2200 189.7250 556.2200 ;
        RECT 196.2400 554.2200 198.2400 556.2200 ;
        RECT 204.7550 554.2200 206.7550 556.2200 ;
        RECT 221.7850 504.5550 223.7850 506.5550 ;
        RECT 213.2700 504.5550 215.2700 506.5550 ;
        RECT 238.8150 497.4600 240.8150 499.4600 ;
        RECT 230.3000 497.4600 232.3000 499.4600 ;
        RECT 221.7850 497.4600 223.7850 499.4600 ;
        RECT 213.2700 497.4600 215.2700 499.4600 ;
        RECT 238.8150 490.3650 240.8150 492.3650 ;
        RECT 230.3000 490.3650 232.3000 492.3650 ;
        RECT 221.7850 490.3650 223.7850 492.3650 ;
        RECT 213.2700 490.3650 215.2700 492.3650 ;
        RECT 230.3000 504.5550 232.3000 506.5550 ;
        RECT 238.8150 504.5550 240.8150 506.5550 ;
        RECT 213.2700 511.6500 215.2700 513.6500 ;
        RECT 221.7850 511.6500 223.7850 513.6500 ;
        RECT 230.3000 511.6500 232.3000 513.6500 ;
        RECT 238.8150 511.6500 240.8150 513.6500 ;
        RECT 213.2700 518.7450 215.2700 520.7450 ;
        RECT 221.7850 518.7450 223.7850 520.7450 ;
        RECT 230.3000 518.7450 232.3000 520.7450 ;
        RECT 238.8150 518.7450 240.8150 520.7450 ;
        RECT 255.8450 504.5550 257.8450 506.5550 ;
        RECT 247.3300 504.5550 249.3300 506.5550 ;
        RECT 272.8750 497.4600 274.8750 499.4600 ;
        RECT 264.3600 497.4600 266.3600 499.4600 ;
        RECT 255.8450 497.4600 257.8450 499.4600 ;
        RECT 247.3300 497.4600 249.3300 499.4600 ;
        RECT 272.8750 490.3650 274.8750 492.3650 ;
        RECT 264.3600 490.3650 266.3600 492.3650 ;
        RECT 255.8450 490.3650 257.8450 492.3650 ;
        RECT 247.3300 490.3650 249.3300 492.3650 ;
        RECT 264.3600 504.5550 266.3600 506.5550 ;
        RECT 272.8750 504.5550 274.8750 506.5550 ;
        RECT 247.3300 511.6500 249.3300 513.6500 ;
        RECT 255.8450 511.6500 257.8450 513.6500 ;
        RECT 264.3600 511.6500 266.3600 513.6500 ;
        RECT 272.8750 511.6500 274.8750 513.6500 ;
        RECT 247.3300 518.7450 249.3300 520.7450 ;
        RECT 255.8450 518.7450 257.8450 520.7450 ;
        RECT 264.3600 518.7450 266.3600 520.7450 ;
        RECT 272.8750 518.7450 274.8750 520.7450 ;
        RECT 221.7850 540.0300 223.7850 542.0300 ;
        RECT 213.2700 540.0300 215.2700 542.0300 ;
        RECT 238.8150 532.9350 240.8150 534.9350 ;
        RECT 230.3000 532.9350 232.3000 534.9350 ;
        RECT 221.7850 532.9350 223.7850 534.9350 ;
        RECT 213.2700 532.9350 215.2700 534.9350 ;
        RECT 238.8150 525.8400 240.8150 527.8400 ;
        RECT 230.3000 525.8400 232.3000 527.8400 ;
        RECT 221.7850 525.8400 223.7850 527.8400 ;
        RECT 213.2700 525.8400 215.2700 527.8400 ;
        RECT 230.3000 540.0300 232.3000 542.0300 ;
        RECT 238.8150 540.0300 240.8150 542.0300 ;
        RECT 213.2700 547.1250 215.2700 549.1250 ;
        RECT 221.7850 547.1250 223.7850 549.1250 ;
        RECT 230.3000 547.1250 232.3000 549.1250 ;
        RECT 238.8150 547.1250 240.8150 549.1250 ;
        RECT 213.2700 554.2200 215.2700 556.2200 ;
        RECT 221.7850 554.2200 223.7850 556.2200 ;
        RECT 230.3000 554.2200 232.3000 556.2200 ;
        RECT 238.8150 554.2200 240.8150 556.2200 ;
        RECT 255.8450 540.0300 257.8450 542.0300 ;
        RECT 247.3300 540.0300 249.3300 542.0300 ;
        RECT 272.8750 532.9350 274.8750 534.9350 ;
        RECT 264.3600 532.9350 266.3600 534.9350 ;
        RECT 255.8450 532.9350 257.8450 534.9350 ;
        RECT 247.3300 532.9350 249.3300 534.9350 ;
        RECT 272.8750 525.8400 274.8750 527.8400 ;
        RECT 264.3600 525.8400 266.3600 527.8400 ;
        RECT 255.8450 525.8400 257.8450 527.8400 ;
        RECT 247.3300 525.8400 249.3300 527.8400 ;
        RECT 264.3600 540.0300 266.3600 542.0300 ;
        RECT 272.8750 540.0300 274.8750 542.0300 ;
        RECT 247.3300 547.1250 249.3300 549.1250 ;
        RECT 255.8450 547.1250 257.8450 549.1250 ;
        RECT 264.3600 547.1250 266.3600 549.1250 ;
        RECT 272.8750 547.1250 274.8750 549.1250 ;
        RECT 247.3300 554.2200 249.3300 556.2200 ;
        RECT 255.8450 554.2200 257.8450 556.2200 ;
        RECT 264.3600 554.2200 266.3600 556.2200 ;
        RECT 272.8750 554.2200 274.8750 556.2200 ;
        RECT 344.0000 419.4150 346.0000 421.4150 ;
        RECT 394.0000 419.4150 396.0000 421.4150 ;
        RECT 281.3900 419.4150 283.3900 421.4150 ;
        RECT 289.9050 419.4150 291.9050 421.4150 ;
        RECT 298.4200 419.4150 300.4200 421.4150 ;
        RECT 306.9350 419.4150 308.9350 421.4150 ;
        RECT 315.4500 419.4150 317.4500 421.4150 ;
        RECT 323.9650 419.4150 325.9650 421.4150 ;
        RECT 414.1500 419.4150 416.1500 421.4150 ;
        RECT 487.5000 419.4150 489.5000 421.4150 ;
        RECT 479.3500 419.4150 481.3500 421.4150 ;
        RECT 471.2000 419.4150 473.2000 421.4150 ;
        RECT 463.0500 419.4150 465.0500 421.4150 ;
        RECT 454.9000 419.4150 456.9000 421.4150 ;
        RECT 446.7500 419.4150 448.7500 421.4150 ;
        RECT 438.6000 419.4150 440.6000 421.4150 ;
        RECT 430.4500 419.4150 432.4500 421.4150 ;
        RECT 422.3000 419.4150 424.3000 421.4150 ;
        RECT 520.1000 419.4150 522.1000 421.4150 ;
        RECT 511.9500 419.4150 513.9500 421.4150 ;
        RECT 503.8000 419.4150 505.8000 421.4150 ;
        RECT 495.6500 419.4150 497.6500 421.4150 ;
        RECT 528.2500 419.4150 530.2500 421.4150 ;
        RECT 536.4000 419.4150 538.4000 421.4150 ;
        RECT 544.5500 419.4150 546.5500 421.4150 ;
        RECT 552.7000 419.4150 554.7000 421.4150 ;
        RECT 394.0000 348.4650 396.0000 350.4650 ;
        RECT 414.1500 348.4650 416.1500 350.4650 ;
        RECT 306.9350 291.7050 308.9350 293.7050 ;
        RECT 298.4200 291.7050 300.4200 293.7050 ;
        RECT 289.9050 291.7050 291.9050 293.7050 ;
        RECT 281.3900 291.7050 283.3900 293.7050 ;
        RECT 306.9350 284.6100 308.9350 286.6100 ;
        RECT 298.4200 284.6100 300.4200 286.6100 ;
        RECT 289.9050 284.6100 291.9050 286.6100 ;
        RECT 281.3900 284.6100 283.3900 286.6100 ;
        RECT 289.9050 298.8000 291.9050 300.8000 ;
        RECT 281.3900 298.8000 283.3900 300.8000 ;
        RECT 298.4200 298.8000 300.4200 300.8000 ;
        RECT 306.9350 298.8000 308.9350 300.8000 ;
        RECT 281.3900 305.8950 283.3900 307.8950 ;
        RECT 289.9050 305.8950 291.9050 307.8950 ;
        RECT 298.4200 305.8950 300.4200 307.8950 ;
        RECT 306.9350 305.8950 308.9350 307.8950 ;
        RECT 281.3900 312.9900 283.3900 314.9900 ;
        RECT 289.9050 312.9900 291.9050 314.9900 ;
        RECT 298.4200 312.9900 300.4200 314.9900 ;
        RECT 306.9350 312.9900 308.9350 314.9900 ;
        RECT 323.9650 291.7050 325.9650 293.7050 ;
        RECT 315.4500 291.7050 317.4500 293.7050 ;
        RECT 323.9650 284.6100 325.9650 286.6100 ;
        RECT 315.4500 284.6100 317.4500 286.6100 ;
        RECT 344.0000 291.7050 346.0000 293.7050 ;
        RECT 344.0000 284.6100 346.0000 286.6100 ;
        RECT 315.4500 298.8000 317.4500 300.8000 ;
        RECT 323.9650 298.8000 325.9650 300.8000 ;
        RECT 315.4500 305.8950 317.4500 307.8950 ;
        RECT 323.9650 305.8950 325.9650 307.8950 ;
        RECT 315.4500 312.9900 317.4500 314.9900 ;
        RECT 323.9650 312.9900 325.9650 314.9900 ;
        RECT 344.0000 312.9900 346.0000 314.9900 ;
        RECT 344.0000 305.8950 346.0000 307.8950 ;
        RECT 344.0000 298.8000 346.0000 300.8000 ;
        RECT 281.3900 320.0850 283.3900 322.0850 ;
        RECT 289.9050 320.0850 291.9050 322.0850 ;
        RECT 298.4200 320.0850 300.4200 322.0850 ;
        RECT 306.9350 320.0850 308.9350 322.0850 ;
        RECT 281.3900 327.1800 283.3900 329.1800 ;
        RECT 289.9050 327.1800 291.9050 329.1800 ;
        RECT 298.4200 327.1800 300.4200 329.1800 ;
        RECT 306.9350 327.1800 308.9350 329.1800 ;
        RECT 323.9650 327.1800 325.9650 329.1800 ;
        RECT 315.4500 327.1800 317.4500 329.1800 ;
        RECT 323.9650 320.0850 325.9650 322.0850 ;
        RECT 315.4500 320.0850 317.4500 322.0850 ;
        RECT 344.0000 327.1800 346.0000 329.1800 ;
        RECT 344.0000 320.0850 346.0000 322.0850 ;
        RECT 344.0000 334.2750 346.0000 336.2750 ;
        RECT 344.0000 341.3700 346.0000 343.3700 ;
        RECT 394.0000 284.6100 396.0000 286.6100 ;
        RECT 394.0000 291.7050 396.0000 293.7050 ;
        RECT 414.1500 284.6100 416.1500 286.6100 ;
        RECT 414.1500 291.7050 416.1500 293.7050 ;
        RECT 394.0000 312.9900 396.0000 314.9900 ;
        RECT 394.0000 305.8950 396.0000 307.8950 ;
        RECT 394.0000 298.8000 396.0000 300.8000 ;
        RECT 414.1500 298.8000 416.1500 300.8000 ;
        RECT 414.1500 305.8950 416.1500 307.8950 ;
        RECT 414.1500 312.9900 416.1500 314.9900 ;
        RECT 394.0000 327.1800 396.0000 329.1800 ;
        RECT 394.0000 320.0850 396.0000 322.0850 ;
        RECT 414.1500 327.1800 416.1500 329.1800 ;
        RECT 414.1500 320.0850 416.1500 322.0850 ;
        RECT 394.0000 334.2750 396.0000 336.2750 ;
        RECT 394.0000 341.3700 396.0000 343.3700 ;
        RECT 414.1500 334.2750 416.1500 336.2750 ;
        RECT 414.1500 341.3700 416.1500 343.3700 ;
        RECT 281.3900 412.3200 283.3900 414.3200 ;
        RECT 289.9050 412.3200 291.9050 414.3200 ;
        RECT 298.4200 412.3200 300.4200 414.3200 ;
        RECT 306.9350 412.3200 308.9350 414.3200 ;
        RECT 344.0000 398.1300 346.0000 400.1300 ;
        RECT 344.0000 412.3200 346.0000 414.3200 ;
        RECT 344.0000 405.2250 346.0000 407.2250 ;
        RECT 315.4500 412.3200 317.4500 414.3200 ;
        RECT 323.9650 412.3200 325.9650 414.3200 ;
        RECT 394.0000 383.9400 396.0000 385.9400 ;
        RECT 414.1500 383.9400 416.1500 385.9400 ;
        RECT 394.0000 355.5600 396.0000 357.5600 ;
        RECT 394.0000 362.6550 396.0000 364.6550 ;
        RECT 414.1500 362.6550 416.1500 364.6550 ;
        RECT 414.1500 355.5600 416.1500 357.5600 ;
        RECT 394.0000 369.7500 396.0000 371.7500 ;
        RECT 394.0000 376.8450 396.0000 378.8450 ;
        RECT 414.1500 376.8450 416.1500 378.8450 ;
        RECT 414.1500 369.7500 416.1500 371.7500 ;
        RECT 394.0000 391.0350 396.0000 393.0350 ;
        RECT 394.0000 398.1300 396.0000 400.1300 ;
        RECT 414.1500 391.0350 416.1500 393.0350 ;
        RECT 414.1500 398.1300 416.1500 400.1300 ;
        RECT 394.0000 405.2250 396.0000 407.2250 ;
        RECT 394.0000 412.3200 396.0000 414.3200 ;
        RECT 414.1500 405.2250 416.1500 407.2250 ;
        RECT 414.1500 412.3200 416.1500 414.3200 ;
        RECT 487.5000 348.4650 489.5000 350.4650 ;
        RECT 479.3500 348.4650 481.3500 350.4650 ;
        RECT 471.2000 348.4650 473.2000 350.4650 ;
        RECT 463.0500 348.4650 465.0500 350.4650 ;
        RECT 454.9000 348.4650 456.9000 350.4650 ;
        RECT 446.7500 348.4650 448.7500 350.4650 ;
        RECT 438.6000 348.4650 440.6000 350.4650 ;
        RECT 430.4500 348.4650 432.4500 350.4650 ;
        RECT 422.3000 348.4650 424.3000 350.4650 ;
        RECT 520.1000 348.4650 522.1000 350.4650 ;
        RECT 511.9500 348.4650 513.9500 350.4650 ;
        RECT 503.8000 348.4650 505.8000 350.4650 ;
        RECT 495.6500 348.4650 497.6500 350.4650 ;
        RECT 528.2500 348.4650 530.2500 350.4650 ;
        RECT 536.4000 348.4650 538.4000 350.4650 ;
        RECT 544.5500 348.4650 546.5500 350.4650 ;
        RECT 552.7000 348.4650 554.7000 350.4650 ;
        RECT 454.9000 284.6100 456.9000 286.6100 ;
        RECT 454.9000 291.7050 456.9000 293.7050 ;
        RECT 454.9000 298.8000 456.9000 300.8000 ;
        RECT 454.9000 305.8950 456.9000 307.8950 ;
        RECT 454.9000 312.9900 456.9000 314.9900 ;
        RECT 446.7500 291.7050 448.7500 293.7050 ;
        RECT 438.6000 291.7050 440.6000 293.7050 ;
        RECT 430.4500 291.7050 432.4500 293.7050 ;
        RECT 422.3000 291.7050 424.3000 293.7050 ;
        RECT 446.7500 284.6100 448.7500 286.6100 ;
        RECT 438.6000 284.6100 440.6000 286.6100 ;
        RECT 430.4500 284.6100 432.4500 286.6100 ;
        RECT 422.3000 284.6100 424.3000 286.6100 ;
        RECT 430.4500 298.8000 432.4500 300.8000 ;
        RECT 422.3000 298.8000 424.3000 300.8000 ;
        RECT 438.6000 298.8000 440.6000 300.8000 ;
        RECT 446.7500 298.8000 448.7500 300.8000 ;
        RECT 422.3000 305.8950 424.3000 307.8950 ;
        RECT 430.4500 305.8950 432.4500 307.8950 ;
        RECT 438.6000 305.8950 440.6000 307.8950 ;
        RECT 446.7500 305.8950 448.7500 307.8950 ;
        RECT 422.3000 312.9900 424.3000 314.9900 ;
        RECT 430.4500 312.9900 432.4500 314.9900 ;
        RECT 438.6000 312.9900 440.6000 314.9900 ;
        RECT 446.7500 312.9900 448.7500 314.9900 ;
        RECT 487.5000 291.7050 489.5000 293.7050 ;
        RECT 479.3500 291.7050 481.3500 293.7050 ;
        RECT 471.2000 291.7050 473.2000 293.7050 ;
        RECT 463.0500 291.7050 465.0500 293.7050 ;
        RECT 487.5000 284.6100 489.5000 286.6100 ;
        RECT 479.3500 284.6100 481.3500 286.6100 ;
        RECT 471.2000 284.6100 473.2000 286.6100 ;
        RECT 463.0500 284.6100 465.0500 286.6100 ;
        RECT 471.2000 298.8000 473.2000 300.8000 ;
        RECT 463.0500 298.8000 465.0500 300.8000 ;
        RECT 479.3500 298.8000 481.3500 300.8000 ;
        RECT 487.5000 298.8000 489.5000 300.8000 ;
        RECT 463.0500 305.8950 465.0500 307.8950 ;
        RECT 471.2000 305.8950 473.2000 307.8950 ;
        RECT 479.3500 305.8950 481.3500 307.8950 ;
        RECT 487.5000 305.8950 489.5000 307.8950 ;
        RECT 463.0500 312.9900 465.0500 314.9900 ;
        RECT 471.2000 312.9900 473.2000 314.9900 ;
        RECT 479.3500 312.9900 481.3500 314.9900 ;
        RECT 487.5000 312.9900 489.5000 314.9900 ;
        RECT 454.9000 320.0850 456.9000 322.0850 ;
        RECT 454.9000 327.1800 456.9000 329.1800 ;
        RECT 454.9000 334.2750 456.9000 336.2750 ;
        RECT 454.9000 341.3700 456.9000 343.3700 ;
        RECT 446.7500 327.1800 448.7500 329.1800 ;
        RECT 438.6000 327.1800 440.6000 329.1800 ;
        RECT 430.4500 327.1800 432.4500 329.1800 ;
        RECT 422.3000 327.1800 424.3000 329.1800 ;
        RECT 446.7500 320.0850 448.7500 322.0850 ;
        RECT 438.6000 320.0850 440.6000 322.0850 ;
        RECT 430.4500 320.0850 432.4500 322.0850 ;
        RECT 422.3000 320.0850 424.3000 322.0850 ;
        RECT 430.4500 341.3700 432.4500 343.3700 ;
        RECT 422.3000 341.3700 424.3000 343.3700 ;
        RECT 446.7500 334.2750 448.7500 336.2750 ;
        RECT 438.6000 334.2750 440.6000 336.2750 ;
        RECT 430.4500 334.2750 432.4500 336.2750 ;
        RECT 422.3000 334.2750 424.3000 336.2750 ;
        RECT 438.6000 341.3700 440.6000 343.3700 ;
        RECT 446.7500 341.3700 448.7500 343.3700 ;
        RECT 487.5000 327.1800 489.5000 329.1800 ;
        RECT 479.3500 327.1800 481.3500 329.1800 ;
        RECT 471.2000 327.1800 473.2000 329.1800 ;
        RECT 463.0500 327.1800 465.0500 329.1800 ;
        RECT 487.5000 320.0850 489.5000 322.0850 ;
        RECT 479.3500 320.0850 481.3500 322.0850 ;
        RECT 471.2000 320.0850 473.2000 322.0850 ;
        RECT 463.0500 320.0850 465.0500 322.0850 ;
        RECT 471.2000 341.3700 473.2000 343.3700 ;
        RECT 463.0500 341.3700 465.0500 343.3700 ;
        RECT 487.5000 334.2750 489.5000 336.2750 ;
        RECT 479.3500 334.2750 481.3500 336.2750 ;
        RECT 471.2000 334.2750 473.2000 336.2750 ;
        RECT 463.0500 334.2750 465.0500 336.2750 ;
        RECT 479.3500 341.3700 481.3500 343.3700 ;
        RECT 487.5000 341.3700 489.5000 343.3700 ;
        RECT 520.1000 291.7050 522.1000 293.7050 ;
        RECT 511.9500 291.7050 513.9500 293.7050 ;
        RECT 503.8000 291.7050 505.8000 293.7050 ;
        RECT 495.6500 291.7050 497.6500 293.7050 ;
        RECT 520.1000 284.6100 522.1000 286.6100 ;
        RECT 511.9500 284.6100 513.9500 286.6100 ;
        RECT 503.8000 284.6100 505.8000 286.6100 ;
        RECT 495.6500 284.6100 497.6500 286.6100 ;
        RECT 503.8000 298.8000 505.8000 300.8000 ;
        RECT 495.6500 298.8000 497.6500 300.8000 ;
        RECT 511.9500 298.8000 513.9500 300.8000 ;
        RECT 520.1000 298.8000 522.1000 300.8000 ;
        RECT 495.6500 305.8950 497.6500 307.8950 ;
        RECT 503.8000 305.8950 505.8000 307.8950 ;
        RECT 511.9500 305.8950 513.9500 307.8950 ;
        RECT 520.1000 305.8950 522.1000 307.8950 ;
        RECT 495.6500 312.9900 497.6500 314.9900 ;
        RECT 503.8000 312.9900 505.8000 314.9900 ;
        RECT 511.9500 312.9900 513.9500 314.9900 ;
        RECT 520.1000 312.9900 522.1000 314.9900 ;
        RECT 552.7000 291.7050 554.7000 293.7050 ;
        RECT 544.5500 291.7050 546.5500 293.7050 ;
        RECT 536.4000 291.7050 538.4000 293.7050 ;
        RECT 528.2500 291.7050 530.2500 293.7050 ;
        RECT 552.7000 284.6100 554.7000 286.6100 ;
        RECT 544.5500 284.6100 546.5500 286.6100 ;
        RECT 536.4000 284.6100 538.4000 286.6100 ;
        RECT 528.2500 284.6100 530.2500 286.6100 ;
        RECT 536.4000 298.8000 538.4000 300.8000 ;
        RECT 528.2500 298.8000 530.2500 300.8000 ;
        RECT 544.5500 298.8000 546.5500 300.8000 ;
        RECT 552.7000 298.8000 554.7000 300.8000 ;
        RECT 528.2500 305.8950 530.2500 307.8950 ;
        RECT 536.4000 305.8950 538.4000 307.8950 ;
        RECT 544.5500 305.8950 546.5500 307.8950 ;
        RECT 552.7000 305.8950 554.7000 307.8950 ;
        RECT 528.2500 312.9900 530.2500 314.9900 ;
        RECT 536.4000 312.9900 538.4000 314.9900 ;
        RECT 544.5500 312.9900 546.5500 314.9900 ;
        RECT 552.7000 312.9900 554.7000 314.9900 ;
        RECT 520.1000 327.1800 522.1000 329.1800 ;
        RECT 511.9500 327.1800 513.9500 329.1800 ;
        RECT 503.8000 327.1800 505.8000 329.1800 ;
        RECT 495.6500 327.1800 497.6500 329.1800 ;
        RECT 520.1000 320.0850 522.1000 322.0850 ;
        RECT 511.9500 320.0850 513.9500 322.0850 ;
        RECT 503.8000 320.0850 505.8000 322.0850 ;
        RECT 495.6500 320.0850 497.6500 322.0850 ;
        RECT 503.8000 341.3700 505.8000 343.3700 ;
        RECT 495.6500 341.3700 497.6500 343.3700 ;
        RECT 520.1000 334.2750 522.1000 336.2750 ;
        RECT 511.9500 334.2750 513.9500 336.2750 ;
        RECT 503.8000 334.2750 505.8000 336.2750 ;
        RECT 495.6500 334.2750 497.6500 336.2750 ;
        RECT 511.9500 341.3700 513.9500 343.3700 ;
        RECT 520.1000 341.3700 522.1000 343.3700 ;
        RECT 552.7000 327.1800 554.7000 329.1800 ;
        RECT 544.5500 327.1800 546.5500 329.1800 ;
        RECT 536.4000 327.1800 538.4000 329.1800 ;
        RECT 528.2500 327.1800 530.2500 329.1800 ;
        RECT 552.7000 320.0850 554.7000 322.0850 ;
        RECT 544.5500 320.0850 546.5500 322.0850 ;
        RECT 536.4000 320.0850 538.4000 322.0850 ;
        RECT 528.2500 320.0850 530.2500 322.0850 ;
        RECT 536.4000 341.3700 538.4000 343.3700 ;
        RECT 528.2500 341.3700 530.2500 343.3700 ;
        RECT 552.7000 334.2750 554.7000 336.2750 ;
        RECT 544.5500 334.2750 546.5500 336.2750 ;
        RECT 536.4000 334.2750 538.4000 336.2750 ;
        RECT 528.2500 334.2750 530.2500 336.2750 ;
        RECT 544.5500 341.3700 546.5500 343.3700 ;
        RECT 552.7000 341.3700 554.7000 343.3700 ;
        RECT 422.3000 383.9400 424.3000 385.9400 ;
        RECT 430.4500 383.9400 432.4500 385.9400 ;
        RECT 438.6000 383.9400 440.6000 385.9400 ;
        RECT 446.7500 383.9400 448.7500 385.9400 ;
        RECT 454.9000 383.9400 456.9000 385.9400 ;
        RECT 463.0500 383.9400 465.0500 385.9400 ;
        RECT 471.2000 383.9400 473.2000 385.9400 ;
        RECT 479.3500 383.9400 481.3500 385.9400 ;
        RECT 487.5000 383.9400 489.5000 385.9400 ;
        RECT 454.9000 355.5600 456.9000 357.5600 ;
        RECT 454.9000 362.6550 456.9000 364.6550 ;
        RECT 454.9000 369.7500 456.9000 371.7500 ;
        RECT 454.9000 376.8450 456.9000 378.8450 ;
        RECT 446.7500 362.6550 448.7500 364.6550 ;
        RECT 438.6000 362.6550 440.6000 364.6550 ;
        RECT 430.4500 362.6550 432.4500 364.6550 ;
        RECT 422.3000 362.6550 424.3000 364.6550 ;
        RECT 446.7500 355.5600 448.7500 357.5600 ;
        RECT 438.6000 355.5600 440.6000 357.5600 ;
        RECT 430.4500 355.5600 432.4500 357.5600 ;
        RECT 422.3000 355.5600 424.3000 357.5600 ;
        RECT 430.4500 376.8450 432.4500 378.8450 ;
        RECT 422.3000 376.8450 424.3000 378.8450 ;
        RECT 446.7500 369.7500 448.7500 371.7500 ;
        RECT 438.6000 369.7500 440.6000 371.7500 ;
        RECT 430.4500 369.7500 432.4500 371.7500 ;
        RECT 422.3000 369.7500 424.3000 371.7500 ;
        RECT 438.6000 376.8450 440.6000 378.8450 ;
        RECT 446.7500 376.8450 448.7500 378.8450 ;
        RECT 487.5000 362.6550 489.5000 364.6550 ;
        RECT 479.3500 362.6550 481.3500 364.6550 ;
        RECT 471.2000 362.6550 473.2000 364.6550 ;
        RECT 463.0500 362.6550 465.0500 364.6550 ;
        RECT 487.5000 355.5600 489.5000 357.5600 ;
        RECT 479.3500 355.5600 481.3500 357.5600 ;
        RECT 471.2000 355.5600 473.2000 357.5600 ;
        RECT 463.0500 355.5600 465.0500 357.5600 ;
        RECT 471.2000 376.8450 473.2000 378.8450 ;
        RECT 463.0500 376.8450 465.0500 378.8450 ;
        RECT 487.5000 369.7500 489.5000 371.7500 ;
        RECT 479.3500 369.7500 481.3500 371.7500 ;
        RECT 471.2000 369.7500 473.2000 371.7500 ;
        RECT 463.0500 369.7500 465.0500 371.7500 ;
        RECT 479.3500 376.8450 481.3500 378.8450 ;
        RECT 487.5000 376.8450 489.5000 378.8450 ;
        RECT 454.9000 391.0350 456.9000 393.0350 ;
        RECT 454.9000 398.1300 456.9000 400.1300 ;
        RECT 454.9000 405.2250 456.9000 407.2250 ;
        RECT 454.9000 412.3200 456.9000 414.3200 ;
        RECT 446.7500 398.1300 448.7500 400.1300 ;
        RECT 438.6000 398.1300 440.6000 400.1300 ;
        RECT 430.4500 398.1300 432.4500 400.1300 ;
        RECT 422.3000 398.1300 424.3000 400.1300 ;
        RECT 446.7500 391.0350 448.7500 393.0350 ;
        RECT 438.6000 391.0350 440.6000 393.0350 ;
        RECT 430.4500 391.0350 432.4500 393.0350 ;
        RECT 422.3000 391.0350 424.3000 393.0350 ;
        RECT 430.4500 412.3200 432.4500 414.3200 ;
        RECT 422.3000 412.3200 424.3000 414.3200 ;
        RECT 446.7500 405.2250 448.7500 407.2250 ;
        RECT 438.6000 405.2250 440.6000 407.2250 ;
        RECT 430.4500 405.2250 432.4500 407.2250 ;
        RECT 422.3000 405.2250 424.3000 407.2250 ;
        RECT 438.6000 412.3200 440.6000 414.3200 ;
        RECT 446.7500 412.3200 448.7500 414.3200 ;
        RECT 487.5000 398.1300 489.5000 400.1300 ;
        RECT 479.3500 398.1300 481.3500 400.1300 ;
        RECT 471.2000 398.1300 473.2000 400.1300 ;
        RECT 463.0500 398.1300 465.0500 400.1300 ;
        RECT 487.5000 391.0350 489.5000 393.0350 ;
        RECT 479.3500 391.0350 481.3500 393.0350 ;
        RECT 471.2000 391.0350 473.2000 393.0350 ;
        RECT 463.0500 391.0350 465.0500 393.0350 ;
        RECT 471.2000 412.3200 473.2000 414.3200 ;
        RECT 463.0500 412.3200 465.0500 414.3200 ;
        RECT 487.5000 405.2250 489.5000 407.2250 ;
        RECT 479.3500 405.2250 481.3500 407.2250 ;
        RECT 471.2000 405.2250 473.2000 407.2250 ;
        RECT 463.0500 405.2250 465.0500 407.2250 ;
        RECT 479.3500 412.3200 481.3500 414.3200 ;
        RECT 487.5000 412.3200 489.5000 414.3200 ;
        RECT 495.6500 383.9400 497.6500 385.9400 ;
        RECT 503.8000 383.9400 505.8000 385.9400 ;
        RECT 511.9500 383.9400 513.9500 385.9400 ;
        RECT 520.1000 383.9400 522.1000 385.9400 ;
        RECT 528.2500 383.9400 530.2500 385.9400 ;
        RECT 536.4000 383.9400 538.4000 385.9400 ;
        RECT 544.5500 383.9400 546.5500 385.9400 ;
        RECT 552.7000 383.9400 554.7000 385.9400 ;
        RECT 520.1000 362.6550 522.1000 364.6550 ;
        RECT 511.9500 362.6550 513.9500 364.6550 ;
        RECT 503.8000 362.6550 505.8000 364.6550 ;
        RECT 495.6500 362.6550 497.6500 364.6550 ;
        RECT 520.1000 355.5600 522.1000 357.5600 ;
        RECT 511.9500 355.5600 513.9500 357.5600 ;
        RECT 503.8000 355.5600 505.8000 357.5600 ;
        RECT 495.6500 355.5600 497.6500 357.5600 ;
        RECT 503.8000 376.8450 505.8000 378.8450 ;
        RECT 495.6500 376.8450 497.6500 378.8450 ;
        RECT 520.1000 369.7500 522.1000 371.7500 ;
        RECT 511.9500 369.7500 513.9500 371.7500 ;
        RECT 503.8000 369.7500 505.8000 371.7500 ;
        RECT 495.6500 369.7500 497.6500 371.7500 ;
        RECT 511.9500 376.8450 513.9500 378.8450 ;
        RECT 520.1000 376.8450 522.1000 378.8450 ;
        RECT 552.7000 362.6550 554.7000 364.6550 ;
        RECT 544.5500 362.6550 546.5500 364.6550 ;
        RECT 536.4000 362.6550 538.4000 364.6550 ;
        RECT 528.2500 362.6550 530.2500 364.6550 ;
        RECT 552.7000 355.5600 554.7000 357.5600 ;
        RECT 544.5500 355.5600 546.5500 357.5600 ;
        RECT 536.4000 355.5600 538.4000 357.5600 ;
        RECT 528.2500 355.5600 530.2500 357.5600 ;
        RECT 536.4000 376.8450 538.4000 378.8450 ;
        RECT 528.2500 376.8450 530.2500 378.8450 ;
        RECT 552.7000 369.7500 554.7000 371.7500 ;
        RECT 544.5500 369.7500 546.5500 371.7500 ;
        RECT 536.4000 369.7500 538.4000 371.7500 ;
        RECT 528.2500 369.7500 530.2500 371.7500 ;
        RECT 544.5500 376.8450 546.5500 378.8450 ;
        RECT 552.7000 376.8450 554.7000 378.8450 ;
        RECT 520.1000 398.1300 522.1000 400.1300 ;
        RECT 511.9500 398.1300 513.9500 400.1300 ;
        RECT 503.8000 398.1300 505.8000 400.1300 ;
        RECT 495.6500 398.1300 497.6500 400.1300 ;
        RECT 520.1000 391.0350 522.1000 393.0350 ;
        RECT 511.9500 391.0350 513.9500 393.0350 ;
        RECT 503.8000 391.0350 505.8000 393.0350 ;
        RECT 495.6500 391.0350 497.6500 393.0350 ;
        RECT 503.8000 412.3200 505.8000 414.3200 ;
        RECT 495.6500 412.3200 497.6500 414.3200 ;
        RECT 520.1000 405.2250 522.1000 407.2250 ;
        RECT 511.9500 405.2250 513.9500 407.2250 ;
        RECT 503.8000 405.2250 505.8000 407.2250 ;
        RECT 495.6500 405.2250 497.6500 407.2250 ;
        RECT 511.9500 412.3200 513.9500 414.3200 ;
        RECT 520.1000 412.3200 522.1000 414.3200 ;
        RECT 552.7000 398.1300 554.7000 400.1300 ;
        RECT 544.5500 398.1300 546.5500 400.1300 ;
        RECT 536.4000 398.1300 538.4000 400.1300 ;
        RECT 528.2500 398.1300 530.2500 400.1300 ;
        RECT 552.7000 391.0350 554.7000 393.0350 ;
        RECT 544.5500 391.0350 546.5500 393.0350 ;
        RECT 536.4000 391.0350 538.4000 393.0350 ;
        RECT 528.2500 391.0350 530.2500 393.0350 ;
        RECT 536.4000 412.3200 538.4000 414.3200 ;
        RECT 528.2500 412.3200 530.2500 414.3200 ;
        RECT 552.7000 405.2250 554.7000 407.2250 ;
        RECT 544.5500 405.2250 546.5500 407.2250 ;
        RECT 536.4000 405.2250 538.4000 407.2250 ;
        RECT 528.2500 405.2250 530.2500 407.2250 ;
        RECT 544.5500 412.3200 546.5500 414.3200 ;
        RECT 552.7000 412.3200 554.7000 414.3200 ;
        RECT 344.0000 454.8900 346.0000 456.8900 ;
        RECT 281.3900 454.8900 283.3900 456.8900 ;
        RECT 289.9050 454.8900 291.9050 456.8900 ;
        RECT 298.4200 454.8900 300.4200 456.8900 ;
        RECT 306.9350 454.8900 308.9350 456.8900 ;
        RECT 315.4500 454.8900 317.4500 456.8900 ;
        RECT 323.9650 454.8900 325.9650 456.8900 ;
        RECT 306.9350 433.6050 308.9350 435.6050 ;
        RECT 298.4200 433.6050 300.4200 435.6050 ;
        RECT 289.9050 433.6050 291.9050 435.6050 ;
        RECT 281.3900 433.6050 283.3900 435.6050 ;
        RECT 306.9350 426.5100 308.9350 428.5100 ;
        RECT 298.4200 426.5100 300.4200 428.5100 ;
        RECT 289.9050 426.5100 291.9050 428.5100 ;
        RECT 281.3900 426.5100 283.3900 428.5100 ;
        RECT 289.9050 447.7950 291.9050 449.7950 ;
        RECT 281.3900 447.7950 283.3900 449.7950 ;
        RECT 306.9350 440.7000 308.9350 442.7000 ;
        RECT 298.4200 440.7000 300.4200 442.7000 ;
        RECT 289.9050 440.7000 291.9050 442.7000 ;
        RECT 281.3900 440.7000 283.3900 442.7000 ;
        RECT 298.4200 447.7950 300.4200 449.7950 ;
        RECT 306.9350 447.7950 308.9350 449.7950 ;
        RECT 323.9650 426.5100 325.9650 428.5100 ;
        RECT 315.4500 426.5100 317.4500 428.5100 ;
        RECT 315.4500 433.6050 317.4500 435.6050 ;
        RECT 323.9650 433.6050 325.9650 435.6050 ;
        RECT 344.0000 426.5100 346.0000 428.5100 ;
        RECT 344.0000 433.6050 346.0000 435.6050 ;
        RECT 315.4500 447.7950 317.4500 449.7950 ;
        RECT 323.9650 440.7000 325.9650 442.7000 ;
        RECT 315.4500 440.7000 317.4500 442.7000 ;
        RECT 323.9650 447.7950 325.9650 449.7950 ;
        RECT 344.0000 440.7000 346.0000 442.7000 ;
        RECT 344.0000 447.7950 346.0000 449.7950 ;
        RECT 306.9350 469.0800 308.9350 471.0800 ;
        RECT 298.4200 469.0800 300.4200 471.0800 ;
        RECT 289.9050 469.0800 291.9050 471.0800 ;
        RECT 281.3900 469.0800 283.3900 471.0800 ;
        RECT 306.9350 461.9850 308.9350 463.9850 ;
        RECT 298.4200 461.9850 300.4200 463.9850 ;
        RECT 289.9050 461.9850 291.9050 463.9850 ;
        RECT 281.3900 461.9850 283.3900 463.9850 ;
        RECT 289.9050 483.2700 291.9050 485.2700 ;
        RECT 281.3900 483.2700 283.3900 485.2700 ;
        RECT 306.9350 476.1750 308.9350 478.1750 ;
        RECT 298.4200 476.1750 300.4200 478.1750 ;
        RECT 289.9050 476.1750 291.9050 478.1750 ;
        RECT 281.3900 476.1750 283.3900 478.1750 ;
        RECT 298.4200 483.2700 300.4200 485.2700 ;
        RECT 306.9350 483.2700 308.9350 485.2700 ;
        RECT 315.4500 469.0800 317.4500 471.0800 ;
        RECT 323.9650 461.9850 325.9650 463.9850 ;
        RECT 315.4500 461.9850 317.4500 463.9850 ;
        RECT 323.9650 469.0800 325.9650 471.0800 ;
        RECT 344.0000 461.9850 346.0000 463.9850 ;
        RECT 344.0000 469.0800 346.0000 471.0800 ;
        RECT 323.9650 483.2700 325.9650 485.2700 ;
        RECT 315.4500 483.2700 317.4500 485.2700 ;
        RECT 323.9650 476.1750 325.9650 478.1750 ;
        RECT 315.4500 476.1750 317.4500 478.1750 ;
        RECT 344.0000 476.1750 346.0000 478.1750 ;
        RECT 344.0000 483.2700 346.0000 485.2700 ;
        RECT 394.0000 454.8900 396.0000 456.8900 ;
        RECT 414.1500 454.8900 416.1500 456.8900 ;
        RECT 394.0000 433.6050 396.0000 435.6050 ;
        RECT 394.0000 426.5100 396.0000 428.5100 ;
        RECT 414.1500 433.6050 416.1500 435.6050 ;
        RECT 414.1500 426.5100 416.1500 428.5100 ;
        RECT 394.0000 447.7950 396.0000 449.7950 ;
        RECT 394.0000 440.7000 396.0000 442.7000 ;
        RECT 414.1500 447.7950 416.1500 449.7950 ;
        RECT 414.1500 440.7000 416.1500 442.7000 ;
        RECT 394.0000 461.9850 396.0000 463.9850 ;
        RECT 394.0000 469.0800 396.0000 471.0800 ;
        RECT 414.1500 461.9850 416.1500 463.9850 ;
        RECT 414.1500 469.0800 416.1500 471.0800 ;
        RECT 394.0000 476.1750 396.0000 478.1750 ;
        RECT 394.0000 483.2700 396.0000 485.2700 ;
        RECT 414.1500 476.1750 416.1500 478.1750 ;
        RECT 414.1500 483.2700 416.1500 485.2700 ;
        RECT 289.9050 504.5550 291.9050 506.5550 ;
        RECT 281.3900 504.5550 283.3900 506.5550 ;
        RECT 306.9350 497.4600 308.9350 499.4600 ;
        RECT 298.4200 497.4600 300.4200 499.4600 ;
        RECT 289.9050 497.4600 291.9050 499.4600 ;
        RECT 281.3900 497.4600 283.3900 499.4600 ;
        RECT 306.9350 490.3650 308.9350 492.3650 ;
        RECT 298.4200 490.3650 300.4200 492.3650 ;
        RECT 289.9050 490.3650 291.9050 492.3650 ;
        RECT 281.3900 490.3650 283.3900 492.3650 ;
        RECT 298.4200 504.5550 300.4200 506.5550 ;
        RECT 306.9350 504.5550 308.9350 506.5550 ;
        RECT 281.3900 511.6500 283.3900 513.6500 ;
        RECT 289.9050 511.6500 291.9050 513.6500 ;
        RECT 298.4200 511.6500 300.4200 513.6500 ;
        RECT 306.9350 511.6500 308.9350 513.6500 ;
        RECT 281.3900 518.7450 283.3900 520.7450 ;
        RECT 289.9050 518.7450 291.9050 520.7450 ;
        RECT 298.4200 518.7450 300.4200 520.7450 ;
        RECT 306.9350 518.7450 308.9350 520.7450 ;
        RECT 315.4500 490.3650 317.4500 492.3650 ;
        RECT 323.9650 490.3650 325.9650 492.3650 ;
        RECT 315.4500 497.4600 317.4500 499.4600 ;
        RECT 323.9650 497.4600 325.9650 499.4600 ;
        RECT 315.4500 504.5550 317.4500 506.5550 ;
        RECT 323.9650 504.5550 325.9650 506.5550 ;
        RECT 344.0000 490.3650 346.0000 492.3650 ;
        RECT 344.0000 497.4600 346.0000 499.4600 ;
        RECT 344.0000 504.5550 346.0000 506.5550 ;
        RECT 323.9650 518.7450 325.9650 520.7450 ;
        RECT 315.4500 518.7450 317.4500 520.7450 ;
        RECT 323.9650 511.6500 325.9650 513.6500 ;
        RECT 315.4500 511.6500 317.4500 513.6500 ;
        RECT 344.0000 511.6500 346.0000 513.6500 ;
        RECT 344.0000 518.7450 346.0000 520.7450 ;
        RECT 289.9050 540.0300 291.9050 542.0300 ;
        RECT 281.3900 540.0300 283.3900 542.0300 ;
        RECT 306.9350 532.9350 308.9350 534.9350 ;
        RECT 298.4200 532.9350 300.4200 534.9350 ;
        RECT 289.9050 532.9350 291.9050 534.9350 ;
        RECT 281.3900 532.9350 283.3900 534.9350 ;
        RECT 306.9350 525.8400 308.9350 527.8400 ;
        RECT 298.4200 525.8400 300.4200 527.8400 ;
        RECT 289.9050 525.8400 291.9050 527.8400 ;
        RECT 281.3900 525.8400 283.3900 527.8400 ;
        RECT 298.4200 540.0300 300.4200 542.0300 ;
        RECT 306.9350 540.0300 308.9350 542.0300 ;
        RECT 281.3900 547.1250 283.3900 549.1250 ;
        RECT 289.9050 547.1250 291.9050 549.1250 ;
        RECT 298.4200 547.1250 300.4200 549.1250 ;
        RECT 306.9350 547.1250 308.9350 549.1250 ;
        RECT 281.3900 554.2200 283.3900 556.2200 ;
        RECT 289.9050 554.2200 291.9050 556.2200 ;
        RECT 298.4200 554.2200 300.4200 556.2200 ;
        RECT 306.9350 554.2200 308.9350 556.2200 ;
        RECT 323.9650 525.8400 325.9650 527.8400 ;
        RECT 315.4500 525.8400 317.4500 527.8400 ;
        RECT 315.4500 532.9350 317.4500 534.9350 ;
        RECT 323.9650 532.9350 325.9650 534.9350 ;
        RECT 315.4500 540.0300 317.4500 542.0300 ;
        RECT 323.9650 540.0300 325.9650 542.0300 ;
        RECT 344.0000 525.8400 346.0000 527.8400 ;
        RECT 344.0000 532.9350 346.0000 534.9350 ;
        RECT 344.0000 540.0300 346.0000 542.0300 ;
        RECT 323.9650 554.2200 325.9650 556.2200 ;
        RECT 315.4500 554.2200 317.4500 556.2200 ;
        RECT 323.9650 547.1250 325.9650 549.1250 ;
        RECT 315.4500 547.1250 317.4500 549.1250 ;
        RECT 344.0000 547.1250 346.0000 549.1250 ;
        RECT 344.0000 554.2200 346.0000 556.2200 ;
        RECT 394.0000 504.5550 396.0000 506.5550 ;
        RECT 394.0000 497.4600 396.0000 499.4600 ;
        RECT 394.0000 490.3650 396.0000 492.3650 ;
        RECT 414.1500 490.3650 416.1500 492.3650 ;
        RECT 414.1500 497.4600 416.1500 499.4600 ;
        RECT 414.1500 504.5550 416.1500 506.5550 ;
        RECT 394.0000 518.7450 396.0000 520.7450 ;
        RECT 394.0000 511.6500 396.0000 513.6500 ;
        RECT 414.1500 518.7450 416.1500 520.7450 ;
        RECT 414.1500 511.6500 416.1500 513.6500 ;
        RECT 394.0000 540.0300 396.0000 542.0300 ;
        RECT 394.0000 532.9350 396.0000 534.9350 ;
        RECT 394.0000 525.8400 396.0000 527.8400 ;
        RECT 414.1500 532.9350 416.1500 534.9350 ;
        RECT 414.1500 525.8400 416.1500 527.8400 ;
        RECT 414.1500 540.0300 416.1500 542.0300 ;
        RECT 394.0000 554.2200 396.0000 556.2200 ;
        RECT 394.0000 547.1250 396.0000 549.1250 ;
        RECT 414.1500 554.2200 416.1500 556.2200 ;
        RECT 414.1500 547.1250 416.1500 549.1250 ;
        RECT 422.3000 454.8900 424.3000 456.8900 ;
        RECT 430.4500 454.8900 432.4500 456.8900 ;
        RECT 438.6000 454.8900 440.6000 456.8900 ;
        RECT 446.7500 454.8900 448.7500 456.8900 ;
        RECT 454.9000 454.8900 456.9000 456.8900 ;
        RECT 463.0500 454.8900 465.0500 456.8900 ;
        RECT 471.2000 454.8900 473.2000 456.8900 ;
        RECT 479.3500 454.8900 481.3500 456.8900 ;
        RECT 487.5000 454.8900 489.5000 456.8900 ;
        RECT 454.9000 426.5100 456.9000 428.5100 ;
        RECT 454.9000 433.6050 456.9000 435.6050 ;
        RECT 454.9000 440.7000 456.9000 442.7000 ;
        RECT 454.9000 447.7950 456.9000 449.7950 ;
        RECT 446.7500 433.6050 448.7500 435.6050 ;
        RECT 438.6000 433.6050 440.6000 435.6050 ;
        RECT 430.4500 433.6050 432.4500 435.6050 ;
        RECT 422.3000 433.6050 424.3000 435.6050 ;
        RECT 446.7500 426.5100 448.7500 428.5100 ;
        RECT 438.6000 426.5100 440.6000 428.5100 ;
        RECT 430.4500 426.5100 432.4500 428.5100 ;
        RECT 422.3000 426.5100 424.3000 428.5100 ;
        RECT 430.4500 447.7950 432.4500 449.7950 ;
        RECT 422.3000 447.7950 424.3000 449.7950 ;
        RECT 446.7500 440.7000 448.7500 442.7000 ;
        RECT 438.6000 440.7000 440.6000 442.7000 ;
        RECT 430.4500 440.7000 432.4500 442.7000 ;
        RECT 422.3000 440.7000 424.3000 442.7000 ;
        RECT 438.6000 447.7950 440.6000 449.7950 ;
        RECT 446.7500 447.7950 448.7500 449.7950 ;
        RECT 487.5000 433.6050 489.5000 435.6050 ;
        RECT 479.3500 433.6050 481.3500 435.6050 ;
        RECT 471.2000 433.6050 473.2000 435.6050 ;
        RECT 463.0500 433.6050 465.0500 435.6050 ;
        RECT 487.5000 426.5100 489.5000 428.5100 ;
        RECT 479.3500 426.5100 481.3500 428.5100 ;
        RECT 471.2000 426.5100 473.2000 428.5100 ;
        RECT 463.0500 426.5100 465.0500 428.5100 ;
        RECT 471.2000 447.7950 473.2000 449.7950 ;
        RECT 463.0500 447.7950 465.0500 449.7950 ;
        RECT 487.5000 440.7000 489.5000 442.7000 ;
        RECT 479.3500 440.7000 481.3500 442.7000 ;
        RECT 471.2000 440.7000 473.2000 442.7000 ;
        RECT 463.0500 440.7000 465.0500 442.7000 ;
        RECT 479.3500 447.7950 481.3500 449.7950 ;
        RECT 487.5000 447.7950 489.5000 449.7950 ;
        RECT 454.9000 461.9850 456.9000 463.9850 ;
        RECT 454.9000 469.0800 456.9000 471.0800 ;
        RECT 454.9000 476.1750 456.9000 478.1750 ;
        RECT 454.9000 483.2700 456.9000 485.2700 ;
        RECT 446.7500 469.0800 448.7500 471.0800 ;
        RECT 438.6000 469.0800 440.6000 471.0800 ;
        RECT 430.4500 469.0800 432.4500 471.0800 ;
        RECT 422.3000 469.0800 424.3000 471.0800 ;
        RECT 446.7500 461.9850 448.7500 463.9850 ;
        RECT 438.6000 461.9850 440.6000 463.9850 ;
        RECT 430.4500 461.9850 432.4500 463.9850 ;
        RECT 422.3000 461.9850 424.3000 463.9850 ;
        RECT 430.4500 483.2700 432.4500 485.2700 ;
        RECT 422.3000 483.2700 424.3000 485.2700 ;
        RECT 446.7500 476.1750 448.7500 478.1750 ;
        RECT 438.6000 476.1750 440.6000 478.1750 ;
        RECT 430.4500 476.1750 432.4500 478.1750 ;
        RECT 422.3000 476.1750 424.3000 478.1750 ;
        RECT 438.6000 483.2700 440.6000 485.2700 ;
        RECT 446.7500 483.2700 448.7500 485.2700 ;
        RECT 487.5000 469.0800 489.5000 471.0800 ;
        RECT 479.3500 469.0800 481.3500 471.0800 ;
        RECT 471.2000 469.0800 473.2000 471.0800 ;
        RECT 463.0500 469.0800 465.0500 471.0800 ;
        RECT 487.5000 461.9850 489.5000 463.9850 ;
        RECT 479.3500 461.9850 481.3500 463.9850 ;
        RECT 471.2000 461.9850 473.2000 463.9850 ;
        RECT 463.0500 461.9850 465.0500 463.9850 ;
        RECT 471.2000 483.2700 473.2000 485.2700 ;
        RECT 463.0500 483.2700 465.0500 485.2700 ;
        RECT 487.5000 476.1750 489.5000 478.1750 ;
        RECT 479.3500 476.1750 481.3500 478.1750 ;
        RECT 471.2000 476.1750 473.2000 478.1750 ;
        RECT 463.0500 476.1750 465.0500 478.1750 ;
        RECT 479.3500 483.2700 481.3500 485.2700 ;
        RECT 487.5000 483.2700 489.5000 485.2700 ;
        RECT 495.6500 454.8900 497.6500 456.8900 ;
        RECT 503.8000 454.8900 505.8000 456.8900 ;
        RECT 511.9500 454.8900 513.9500 456.8900 ;
        RECT 520.1000 454.8900 522.1000 456.8900 ;
        RECT 528.2500 454.8900 530.2500 456.8900 ;
        RECT 536.4000 454.8900 538.4000 456.8900 ;
        RECT 544.5500 454.8900 546.5500 456.8900 ;
        RECT 552.7000 454.8900 554.7000 456.8900 ;
        RECT 520.1000 433.6050 522.1000 435.6050 ;
        RECT 511.9500 433.6050 513.9500 435.6050 ;
        RECT 503.8000 433.6050 505.8000 435.6050 ;
        RECT 495.6500 433.6050 497.6500 435.6050 ;
        RECT 520.1000 426.5100 522.1000 428.5100 ;
        RECT 511.9500 426.5100 513.9500 428.5100 ;
        RECT 503.8000 426.5100 505.8000 428.5100 ;
        RECT 495.6500 426.5100 497.6500 428.5100 ;
        RECT 503.8000 447.7950 505.8000 449.7950 ;
        RECT 495.6500 447.7950 497.6500 449.7950 ;
        RECT 520.1000 440.7000 522.1000 442.7000 ;
        RECT 511.9500 440.7000 513.9500 442.7000 ;
        RECT 503.8000 440.7000 505.8000 442.7000 ;
        RECT 495.6500 440.7000 497.6500 442.7000 ;
        RECT 511.9500 447.7950 513.9500 449.7950 ;
        RECT 520.1000 447.7950 522.1000 449.7950 ;
        RECT 552.7000 433.6050 554.7000 435.6050 ;
        RECT 544.5500 433.6050 546.5500 435.6050 ;
        RECT 536.4000 433.6050 538.4000 435.6050 ;
        RECT 528.2500 433.6050 530.2500 435.6050 ;
        RECT 552.7000 426.5100 554.7000 428.5100 ;
        RECT 544.5500 426.5100 546.5500 428.5100 ;
        RECT 536.4000 426.5100 538.4000 428.5100 ;
        RECT 528.2500 426.5100 530.2500 428.5100 ;
        RECT 536.4000 447.7950 538.4000 449.7950 ;
        RECT 528.2500 447.7950 530.2500 449.7950 ;
        RECT 552.7000 440.7000 554.7000 442.7000 ;
        RECT 544.5500 440.7000 546.5500 442.7000 ;
        RECT 536.4000 440.7000 538.4000 442.7000 ;
        RECT 528.2500 440.7000 530.2500 442.7000 ;
        RECT 544.5500 447.7950 546.5500 449.7950 ;
        RECT 552.7000 447.7950 554.7000 449.7950 ;
        RECT 520.1000 469.0800 522.1000 471.0800 ;
        RECT 511.9500 469.0800 513.9500 471.0800 ;
        RECT 503.8000 469.0800 505.8000 471.0800 ;
        RECT 495.6500 469.0800 497.6500 471.0800 ;
        RECT 520.1000 461.9850 522.1000 463.9850 ;
        RECT 511.9500 461.9850 513.9500 463.9850 ;
        RECT 503.8000 461.9850 505.8000 463.9850 ;
        RECT 495.6500 461.9850 497.6500 463.9850 ;
        RECT 503.8000 483.2700 505.8000 485.2700 ;
        RECT 495.6500 483.2700 497.6500 485.2700 ;
        RECT 520.1000 476.1750 522.1000 478.1750 ;
        RECT 511.9500 476.1750 513.9500 478.1750 ;
        RECT 503.8000 476.1750 505.8000 478.1750 ;
        RECT 495.6500 476.1750 497.6500 478.1750 ;
        RECT 511.9500 483.2700 513.9500 485.2700 ;
        RECT 520.1000 483.2700 522.1000 485.2700 ;
        RECT 552.7000 469.0800 554.7000 471.0800 ;
        RECT 544.5500 469.0800 546.5500 471.0800 ;
        RECT 536.4000 469.0800 538.4000 471.0800 ;
        RECT 528.2500 469.0800 530.2500 471.0800 ;
        RECT 552.7000 461.9850 554.7000 463.9850 ;
        RECT 544.5500 461.9850 546.5500 463.9850 ;
        RECT 536.4000 461.9850 538.4000 463.9850 ;
        RECT 528.2500 461.9850 530.2500 463.9850 ;
        RECT 536.4000 483.2700 538.4000 485.2700 ;
        RECT 528.2500 483.2700 530.2500 485.2700 ;
        RECT 552.7000 476.1750 554.7000 478.1750 ;
        RECT 544.5500 476.1750 546.5500 478.1750 ;
        RECT 536.4000 476.1750 538.4000 478.1750 ;
        RECT 528.2500 476.1750 530.2500 478.1750 ;
        RECT 544.5500 483.2700 546.5500 485.2700 ;
        RECT 552.7000 483.2700 554.7000 485.2700 ;
        RECT 454.9000 490.3650 456.9000 492.3650 ;
        RECT 454.9000 497.4600 456.9000 499.4600 ;
        RECT 454.9000 504.5550 456.9000 506.5550 ;
        RECT 454.9000 511.6500 456.9000 513.6500 ;
        RECT 454.9000 518.7450 456.9000 520.7450 ;
        RECT 430.4500 504.5550 432.4500 506.5550 ;
        RECT 422.3000 504.5550 424.3000 506.5550 ;
        RECT 446.7500 497.4600 448.7500 499.4600 ;
        RECT 438.6000 497.4600 440.6000 499.4600 ;
        RECT 430.4500 497.4600 432.4500 499.4600 ;
        RECT 422.3000 497.4600 424.3000 499.4600 ;
        RECT 446.7500 490.3650 448.7500 492.3650 ;
        RECT 438.6000 490.3650 440.6000 492.3650 ;
        RECT 430.4500 490.3650 432.4500 492.3650 ;
        RECT 422.3000 490.3650 424.3000 492.3650 ;
        RECT 438.6000 504.5550 440.6000 506.5550 ;
        RECT 446.7500 504.5550 448.7500 506.5550 ;
        RECT 422.3000 511.6500 424.3000 513.6500 ;
        RECT 430.4500 511.6500 432.4500 513.6500 ;
        RECT 438.6000 511.6500 440.6000 513.6500 ;
        RECT 446.7500 511.6500 448.7500 513.6500 ;
        RECT 422.3000 518.7450 424.3000 520.7450 ;
        RECT 430.4500 518.7450 432.4500 520.7450 ;
        RECT 438.6000 518.7450 440.6000 520.7450 ;
        RECT 446.7500 518.7450 448.7500 520.7450 ;
        RECT 471.2000 504.5550 473.2000 506.5550 ;
        RECT 463.0500 504.5550 465.0500 506.5550 ;
        RECT 487.5000 497.4600 489.5000 499.4600 ;
        RECT 479.3500 497.4600 481.3500 499.4600 ;
        RECT 471.2000 497.4600 473.2000 499.4600 ;
        RECT 463.0500 497.4600 465.0500 499.4600 ;
        RECT 487.5000 490.3650 489.5000 492.3650 ;
        RECT 479.3500 490.3650 481.3500 492.3650 ;
        RECT 471.2000 490.3650 473.2000 492.3650 ;
        RECT 463.0500 490.3650 465.0500 492.3650 ;
        RECT 479.3500 504.5550 481.3500 506.5550 ;
        RECT 487.5000 504.5550 489.5000 506.5550 ;
        RECT 463.0500 511.6500 465.0500 513.6500 ;
        RECT 471.2000 511.6500 473.2000 513.6500 ;
        RECT 479.3500 511.6500 481.3500 513.6500 ;
        RECT 487.5000 511.6500 489.5000 513.6500 ;
        RECT 463.0500 518.7450 465.0500 520.7450 ;
        RECT 471.2000 518.7450 473.2000 520.7450 ;
        RECT 479.3500 518.7450 481.3500 520.7450 ;
        RECT 487.5000 518.7450 489.5000 520.7450 ;
        RECT 454.9000 525.8400 456.9000 527.8400 ;
        RECT 454.9000 532.9350 456.9000 534.9350 ;
        RECT 454.9000 540.0300 456.9000 542.0300 ;
        RECT 454.9000 547.1250 456.9000 549.1250 ;
        RECT 454.9000 554.2200 456.9000 556.2200 ;
        RECT 430.4500 540.0300 432.4500 542.0300 ;
        RECT 422.3000 540.0300 424.3000 542.0300 ;
        RECT 446.7500 532.9350 448.7500 534.9350 ;
        RECT 438.6000 532.9350 440.6000 534.9350 ;
        RECT 430.4500 532.9350 432.4500 534.9350 ;
        RECT 422.3000 532.9350 424.3000 534.9350 ;
        RECT 446.7500 525.8400 448.7500 527.8400 ;
        RECT 438.6000 525.8400 440.6000 527.8400 ;
        RECT 430.4500 525.8400 432.4500 527.8400 ;
        RECT 422.3000 525.8400 424.3000 527.8400 ;
        RECT 438.6000 540.0300 440.6000 542.0300 ;
        RECT 446.7500 540.0300 448.7500 542.0300 ;
        RECT 422.3000 547.1250 424.3000 549.1250 ;
        RECT 430.4500 547.1250 432.4500 549.1250 ;
        RECT 438.6000 547.1250 440.6000 549.1250 ;
        RECT 446.7500 547.1250 448.7500 549.1250 ;
        RECT 422.3000 554.2200 424.3000 556.2200 ;
        RECT 430.4500 554.2200 432.4500 556.2200 ;
        RECT 438.6000 554.2200 440.6000 556.2200 ;
        RECT 446.7500 554.2200 448.7500 556.2200 ;
        RECT 471.2000 540.0300 473.2000 542.0300 ;
        RECT 463.0500 540.0300 465.0500 542.0300 ;
        RECT 487.5000 532.9350 489.5000 534.9350 ;
        RECT 479.3500 532.9350 481.3500 534.9350 ;
        RECT 471.2000 532.9350 473.2000 534.9350 ;
        RECT 463.0500 532.9350 465.0500 534.9350 ;
        RECT 487.5000 525.8400 489.5000 527.8400 ;
        RECT 479.3500 525.8400 481.3500 527.8400 ;
        RECT 471.2000 525.8400 473.2000 527.8400 ;
        RECT 463.0500 525.8400 465.0500 527.8400 ;
        RECT 479.3500 540.0300 481.3500 542.0300 ;
        RECT 487.5000 540.0300 489.5000 542.0300 ;
        RECT 463.0500 547.1250 465.0500 549.1250 ;
        RECT 471.2000 547.1250 473.2000 549.1250 ;
        RECT 479.3500 547.1250 481.3500 549.1250 ;
        RECT 487.5000 547.1250 489.5000 549.1250 ;
        RECT 463.0500 554.2200 465.0500 556.2200 ;
        RECT 471.2000 554.2200 473.2000 556.2200 ;
        RECT 479.3500 554.2200 481.3500 556.2200 ;
        RECT 487.5000 554.2200 489.5000 556.2200 ;
        RECT 503.8000 504.5550 505.8000 506.5550 ;
        RECT 495.6500 504.5550 497.6500 506.5550 ;
        RECT 520.1000 497.4600 522.1000 499.4600 ;
        RECT 511.9500 497.4600 513.9500 499.4600 ;
        RECT 503.8000 497.4600 505.8000 499.4600 ;
        RECT 495.6500 497.4600 497.6500 499.4600 ;
        RECT 520.1000 490.3650 522.1000 492.3650 ;
        RECT 511.9500 490.3650 513.9500 492.3650 ;
        RECT 503.8000 490.3650 505.8000 492.3650 ;
        RECT 495.6500 490.3650 497.6500 492.3650 ;
        RECT 511.9500 504.5550 513.9500 506.5550 ;
        RECT 520.1000 504.5550 522.1000 506.5550 ;
        RECT 495.6500 511.6500 497.6500 513.6500 ;
        RECT 503.8000 511.6500 505.8000 513.6500 ;
        RECT 511.9500 511.6500 513.9500 513.6500 ;
        RECT 520.1000 511.6500 522.1000 513.6500 ;
        RECT 495.6500 518.7450 497.6500 520.7450 ;
        RECT 503.8000 518.7450 505.8000 520.7450 ;
        RECT 511.9500 518.7450 513.9500 520.7450 ;
        RECT 520.1000 518.7450 522.1000 520.7450 ;
        RECT 536.4000 504.5550 538.4000 506.5550 ;
        RECT 528.2500 504.5550 530.2500 506.5550 ;
        RECT 552.7000 497.4600 554.7000 499.4600 ;
        RECT 544.5500 497.4600 546.5500 499.4600 ;
        RECT 536.4000 497.4600 538.4000 499.4600 ;
        RECT 528.2500 497.4600 530.2500 499.4600 ;
        RECT 552.7000 490.3650 554.7000 492.3650 ;
        RECT 544.5500 490.3650 546.5500 492.3650 ;
        RECT 536.4000 490.3650 538.4000 492.3650 ;
        RECT 528.2500 490.3650 530.2500 492.3650 ;
        RECT 544.5500 504.5550 546.5500 506.5550 ;
        RECT 552.7000 504.5550 554.7000 506.5550 ;
        RECT 528.2500 511.6500 530.2500 513.6500 ;
        RECT 536.4000 511.6500 538.4000 513.6500 ;
        RECT 544.5500 511.6500 546.5500 513.6500 ;
        RECT 552.7000 511.6500 554.7000 513.6500 ;
        RECT 528.2500 518.7450 530.2500 520.7450 ;
        RECT 536.4000 518.7450 538.4000 520.7450 ;
        RECT 544.5500 518.7450 546.5500 520.7450 ;
        RECT 552.7000 518.7450 554.7000 520.7450 ;
        RECT 503.8000 540.0300 505.8000 542.0300 ;
        RECT 495.6500 540.0300 497.6500 542.0300 ;
        RECT 520.1000 532.9350 522.1000 534.9350 ;
        RECT 511.9500 532.9350 513.9500 534.9350 ;
        RECT 503.8000 532.9350 505.8000 534.9350 ;
        RECT 495.6500 532.9350 497.6500 534.9350 ;
        RECT 520.1000 525.8400 522.1000 527.8400 ;
        RECT 511.9500 525.8400 513.9500 527.8400 ;
        RECT 503.8000 525.8400 505.8000 527.8400 ;
        RECT 495.6500 525.8400 497.6500 527.8400 ;
        RECT 511.9500 540.0300 513.9500 542.0300 ;
        RECT 520.1000 540.0300 522.1000 542.0300 ;
        RECT 495.6500 547.1250 497.6500 549.1250 ;
        RECT 503.8000 547.1250 505.8000 549.1250 ;
        RECT 511.9500 547.1250 513.9500 549.1250 ;
        RECT 520.1000 547.1250 522.1000 549.1250 ;
        RECT 495.6500 554.2200 497.6500 556.2200 ;
        RECT 503.8000 554.2200 505.8000 556.2200 ;
        RECT 511.9500 554.2200 513.9500 556.2200 ;
        RECT 520.1000 554.2200 522.1000 556.2200 ;
        RECT 536.4000 540.0300 538.4000 542.0300 ;
        RECT 528.2500 540.0300 530.2500 542.0300 ;
        RECT 552.7000 532.9350 554.7000 534.9350 ;
        RECT 544.5500 532.9350 546.5500 534.9350 ;
        RECT 536.4000 532.9350 538.4000 534.9350 ;
        RECT 528.2500 532.9350 530.2500 534.9350 ;
        RECT 552.7000 525.8400 554.7000 527.8400 ;
        RECT 544.5500 525.8400 546.5500 527.8400 ;
        RECT 536.4000 525.8400 538.4000 527.8400 ;
        RECT 528.2500 525.8400 530.2500 527.8400 ;
        RECT 544.5500 540.0300 546.5500 542.0300 ;
        RECT 552.7000 540.0300 554.7000 542.0300 ;
        RECT 528.2500 547.1250 530.2500 549.1250 ;
        RECT 536.4000 547.1250 538.4000 549.1250 ;
        RECT 544.5500 547.1250 546.5500 549.1250 ;
        RECT 552.7000 547.1250 554.7000 549.1250 ;
        RECT 528.2500 554.2200 530.2500 556.2200 ;
        RECT 536.4000 554.2200 538.4000 556.2200 ;
        RECT 544.5500 554.2200 546.5500 556.2200 ;
        RECT 552.7000 554.2200 554.7000 556.2200 ;
        RECT 699.4000 64.6650 701.4000 66.6650 ;
        RECT 699.4000 71.7600 701.4000 73.7600 ;
        RECT 699.4000 78.8550 701.4000 80.8550 ;
        RECT 699.4000 85.9500 701.4000 87.9500 ;
        RECT 699.4000 93.0450 701.4000 95.0450 ;
        RECT 699.4000 100.1400 701.4000 102.1400 ;
        RECT 699.4000 107.2350 701.4000 109.2350 ;
        RECT 699.4000 114.3300 701.4000 116.3300 ;
        RECT 699.4000 121.4250 701.4000 123.4250 ;
        RECT 699.4000 128.5200 701.4000 130.5200 ;
        RECT 699.4000 135.6150 701.4000 137.6150 ;
        RECT 626.0500 64.6650 628.0500 66.6650 ;
        RECT 617.9000 64.6650 619.9000 66.6650 ;
        RECT 609.7500 64.6650 611.7500 66.6650 ;
        RECT 601.6000 64.6650 603.6000 66.6650 ;
        RECT 593.4500 64.6650 595.4500 66.6650 ;
        RECT 585.3000 64.6650 587.3000 66.6650 ;
        RECT 577.1500 64.6650 579.1500 66.6650 ;
        RECT 569.0000 64.6650 571.0000 66.6650 ;
        RECT 560.8500 64.6650 562.8500 66.6650 ;
        RECT 658.6500 64.6650 660.6500 66.6650 ;
        RECT 650.5000 64.6650 652.5000 66.6650 ;
        RECT 642.3500 64.6650 644.3500 66.6650 ;
        RECT 634.2000 64.6650 636.2000 66.6650 ;
        RECT 666.8000 64.6650 668.8000 66.6650 ;
        RECT 674.9500 64.6650 676.9500 66.6650 ;
        RECT 683.1000 64.6650 685.1000 66.6650 ;
        RECT 691.2500 64.6650 693.2500 66.6650 ;
        RECT 593.4500 71.7600 595.4500 73.7600 ;
        RECT 593.4500 78.8550 595.4500 80.8550 ;
        RECT 593.4500 85.9500 595.4500 87.9500 ;
        RECT 593.4500 93.0450 595.4500 95.0450 ;
        RECT 593.4500 100.1400 595.4500 102.1400 ;
        RECT 560.8500 85.9500 562.8500 87.9500 ;
        RECT 569.0000 85.9500 571.0000 87.9500 ;
        RECT 577.1500 85.9500 579.1500 87.9500 ;
        RECT 585.3000 85.9500 587.3000 87.9500 ;
        RECT 585.3000 78.8550 587.3000 80.8550 ;
        RECT 577.1500 78.8550 579.1500 80.8550 ;
        RECT 569.0000 78.8550 571.0000 80.8550 ;
        RECT 560.8500 78.8550 562.8500 80.8550 ;
        RECT 585.3000 71.7600 587.3000 73.7600 ;
        RECT 577.1500 71.7600 579.1500 73.7600 ;
        RECT 569.0000 71.7600 571.0000 73.7600 ;
        RECT 560.8500 71.7600 562.8500 73.7600 ;
        RECT 560.8500 93.0450 562.8500 95.0450 ;
        RECT 569.0000 93.0450 571.0000 95.0450 ;
        RECT 577.1500 93.0450 579.1500 95.0450 ;
        RECT 585.3000 93.0450 587.3000 95.0450 ;
        RECT 560.8500 100.1400 562.8500 102.1400 ;
        RECT 569.0000 100.1400 571.0000 102.1400 ;
        RECT 577.1500 100.1400 579.1500 102.1400 ;
        RECT 585.3000 100.1400 587.3000 102.1400 ;
        RECT 601.6000 85.9500 603.6000 87.9500 ;
        RECT 609.7500 85.9500 611.7500 87.9500 ;
        RECT 617.9000 85.9500 619.9000 87.9500 ;
        RECT 626.0500 85.9500 628.0500 87.9500 ;
        RECT 626.0500 78.8550 628.0500 80.8550 ;
        RECT 617.9000 78.8550 619.9000 80.8550 ;
        RECT 609.7500 78.8550 611.7500 80.8550 ;
        RECT 601.6000 78.8550 603.6000 80.8550 ;
        RECT 626.0500 71.7600 628.0500 73.7600 ;
        RECT 617.9000 71.7600 619.9000 73.7600 ;
        RECT 609.7500 71.7600 611.7500 73.7600 ;
        RECT 601.6000 71.7600 603.6000 73.7600 ;
        RECT 601.6000 93.0450 603.6000 95.0450 ;
        RECT 609.7500 93.0450 611.7500 95.0450 ;
        RECT 617.9000 93.0450 619.9000 95.0450 ;
        RECT 626.0500 93.0450 628.0500 95.0450 ;
        RECT 601.6000 100.1400 603.6000 102.1400 ;
        RECT 609.7500 100.1400 611.7500 102.1400 ;
        RECT 617.9000 100.1400 619.9000 102.1400 ;
        RECT 626.0500 100.1400 628.0500 102.1400 ;
        RECT 593.4500 107.2350 595.4500 109.2350 ;
        RECT 593.4500 114.3300 595.4500 116.3300 ;
        RECT 593.4500 121.4250 595.4500 123.4250 ;
        RECT 593.4500 128.5200 595.4500 130.5200 ;
        RECT 593.4500 135.6150 595.4500 137.6150 ;
        RECT 560.8500 121.4250 562.8500 123.4250 ;
        RECT 569.0000 121.4250 571.0000 123.4250 ;
        RECT 577.1500 121.4250 579.1500 123.4250 ;
        RECT 585.3000 121.4250 587.3000 123.4250 ;
        RECT 585.3000 114.3300 587.3000 116.3300 ;
        RECT 577.1500 114.3300 579.1500 116.3300 ;
        RECT 569.0000 114.3300 571.0000 116.3300 ;
        RECT 560.8500 114.3300 562.8500 116.3300 ;
        RECT 585.3000 107.2350 587.3000 109.2350 ;
        RECT 577.1500 107.2350 579.1500 109.2350 ;
        RECT 569.0000 107.2350 571.0000 109.2350 ;
        RECT 560.8500 107.2350 562.8500 109.2350 ;
        RECT 560.8500 128.5200 562.8500 130.5200 ;
        RECT 569.0000 128.5200 571.0000 130.5200 ;
        RECT 577.1500 128.5200 579.1500 130.5200 ;
        RECT 585.3000 128.5200 587.3000 130.5200 ;
        RECT 560.8500 135.6150 562.8500 137.6150 ;
        RECT 569.0000 135.6150 571.0000 137.6150 ;
        RECT 577.1500 135.6150 579.1500 137.6150 ;
        RECT 585.3000 135.6150 587.3000 137.6150 ;
        RECT 601.6000 121.4250 603.6000 123.4250 ;
        RECT 609.7500 121.4250 611.7500 123.4250 ;
        RECT 617.9000 121.4250 619.9000 123.4250 ;
        RECT 626.0500 121.4250 628.0500 123.4250 ;
        RECT 626.0500 114.3300 628.0500 116.3300 ;
        RECT 617.9000 114.3300 619.9000 116.3300 ;
        RECT 609.7500 114.3300 611.7500 116.3300 ;
        RECT 601.6000 114.3300 603.6000 116.3300 ;
        RECT 626.0500 107.2350 628.0500 109.2350 ;
        RECT 617.9000 107.2350 619.9000 109.2350 ;
        RECT 609.7500 107.2350 611.7500 109.2350 ;
        RECT 601.6000 107.2350 603.6000 109.2350 ;
        RECT 601.6000 128.5200 603.6000 130.5200 ;
        RECT 609.7500 128.5200 611.7500 130.5200 ;
        RECT 617.9000 128.5200 619.9000 130.5200 ;
        RECT 626.0500 128.5200 628.0500 130.5200 ;
        RECT 601.6000 135.6150 603.6000 137.6150 ;
        RECT 609.7500 135.6150 611.7500 137.6150 ;
        RECT 617.9000 135.6150 619.9000 137.6150 ;
        RECT 626.0500 135.6150 628.0500 137.6150 ;
        RECT 634.2000 85.9500 636.2000 87.9500 ;
        RECT 642.3500 85.9500 644.3500 87.9500 ;
        RECT 650.5000 85.9500 652.5000 87.9500 ;
        RECT 658.6500 85.9500 660.6500 87.9500 ;
        RECT 658.6500 78.8550 660.6500 80.8550 ;
        RECT 650.5000 78.8550 652.5000 80.8550 ;
        RECT 642.3500 78.8550 644.3500 80.8550 ;
        RECT 634.2000 78.8550 636.2000 80.8550 ;
        RECT 658.6500 71.7600 660.6500 73.7600 ;
        RECT 650.5000 71.7600 652.5000 73.7600 ;
        RECT 642.3500 71.7600 644.3500 73.7600 ;
        RECT 634.2000 71.7600 636.2000 73.7600 ;
        RECT 634.2000 93.0450 636.2000 95.0450 ;
        RECT 642.3500 93.0450 644.3500 95.0450 ;
        RECT 650.5000 93.0450 652.5000 95.0450 ;
        RECT 658.6500 93.0450 660.6500 95.0450 ;
        RECT 634.2000 100.1400 636.2000 102.1400 ;
        RECT 642.3500 100.1400 644.3500 102.1400 ;
        RECT 650.5000 100.1400 652.5000 102.1400 ;
        RECT 658.6500 100.1400 660.6500 102.1400 ;
        RECT 666.8000 85.9500 668.8000 87.9500 ;
        RECT 674.9500 85.9500 676.9500 87.9500 ;
        RECT 683.1000 85.9500 685.1000 87.9500 ;
        RECT 691.2500 85.9500 693.2500 87.9500 ;
        RECT 691.2500 78.8550 693.2500 80.8550 ;
        RECT 683.1000 78.8550 685.1000 80.8550 ;
        RECT 674.9500 78.8550 676.9500 80.8550 ;
        RECT 666.8000 78.8550 668.8000 80.8550 ;
        RECT 691.2500 71.7600 693.2500 73.7600 ;
        RECT 683.1000 71.7600 685.1000 73.7600 ;
        RECT 674.9500 71.7600 676.9500 73.7600 ;
        RECT 666.8000 71.7600 668.8000 73.7600 ;
        RECT 666.8000 93.0450 668.8000 95.0450 ;
        RECT 674.9500 93.0450 676.9500 95.0450 ;
        RECT 683.1000 93.0450 685.1000 95.0450 ;
        RECT 691.2500 93.0450 693.2500 95.0450 ;
        RECT 666.8000 100.1400 668.8000 102.1400 ;
        RECT 674.9500 100.1400 676.9500 102.1400 ;
        RECT 683.1000 100.1400 685.1000 102.1400 ;
        RECT 691.2500 100.1400 693.2500 102.1400 ;
        RECT 634.2000 121.4250 636.2000 123.4250 ;
        RECT 642.3500 121.4250 644.3500 123.4250 ;
        RECT 650.5000 121.4250 652.5000 123.4250 ;
        RECT 658.6500 121.4250 660.6500 123.4250 ;
        RECT 658.6500 114.3300 660.6500 116.3300 ;
        RECT 650.5000 114.3300 652.5000 116.3300 ;
        RECT 642.3500 114.3300 644.3500 116.3300 ;
        RECT 634.2000 114.3300 636.2000 116.3300 ;
        RECT 658.6500 107.2350 660.6500 109.2350 ;
        RECT 650.5000 107.2350 652.5000 109.2350 ;
        RECT 642.3500 107.2350 644.3500 109.2350 ;
        RECT 634.2000 107.2350 636.2000 109.2350 ;
        RECT 634.2000 128.5200 636.2000 130.5200 ;
        RECT 642.3500 128.5200 644.3500 130.5200 ;
        RECT 650.5000 128.5200 652.5000 130.5200 ;
        RECT 658.6500 128.5200 660.6500 130.5200 ;
        RECT 634.2000 135.6150 636.2000 137.6150 ;
        RECT 642.3500 135.6150 644.3500 137.6150 ;
        RECT 650.5000 135.6150 652.5000 137.6150 ;
        RECT 658.6500 135.6150 660.6500 137.6150 ;
        RECT 666.8000 121.4250 668.8000 123.4250 ;
        RECT 674.9500 121.4250 676.9500 123.4250 ;
        RECT 683.1000 121.4250 685.1000 123.4250 ;
        RECT 691.2500 121.4250 693.2500 123.4250 ;
        RECT 691.2500 114.3300 693.2500 116.3300 ;
        RECT 683.1000 114.3300 685.1000 116.3300 ;
        RECT 674.9500 114.3300 676.9500 116.3300 ;
        RECT 666.8000 114.3300 668.8000 116.3300 ;
        RECT 691.2500 107.2350 693.2500 109.2350 ;
        RECT 683.1000 107.2350 685.1000 109.2350 ;
        RECT 674.9500 107.2350 676.9500 109.2350 ;
        RECT 666.8000 107.2350 668.8000 109.2350 ;
        RECT 666.8000 128.5200 668.8000 130.5200 ;
        RECT 674.9500 128.5200 676.9500 130.5200 ;
        RECT 683.1000 128.5200 685.1000 130.5200 ;
        RECT 691.2500 128.5200 693.2500 130.5200 ;
        RECT 666.8000 135.6150 668.8000 137.6150 ;
        RECT 674.9500 135.6150 676.9500 137.6150 ;
        RECT 683.1000 135.6150 685.1000 137.6150 ;
        RECT 691.2500 135.6150 693.2500 137.6150 ;
        RECT 764.6000 64.6650 766.6000 66.6650 ;
        RECT 756.4500 64.6650 758.4500 66.6650 ;
        RECT 748.3000 64.6650 750.3000 66.6650 ;
        RECT 740.1500 64.6650 742.1500 66.6650 ;
        RECT 732.0000 64.6650 734.0000 66.6650 ;
        RECT 723.8500 64.6650 725.8500 66.6650 ;
        RECT 715.7000 64.6650 717.7000 66.6650 ;
        RECT 707.5500 64.6650 709.5500 66.6650 ;
        RECT 805.3500 64.6650 807.3500 66.6650 ;
        RECT 797.2000 64.6650 799.2000 66.6650 ;
        RECT 789.0500 64.6650 791.0500 66.6650 ;
        RECT 780.9000 64.6650 782.9000 66.6650 ;
        RECT 772.7500 64.6650 774.7500 66.6650 ;
        RECT 813.5000 64.6650 815.5000 66.6650 ;
        RECT 821.6500 64.6650 823.6500 66.6650 ;
        RECT 829.8000 64.6650 831.8000 66.6650 ;
        RECT 837.9500 64.6650 839.9500 66.6650 ;
        RECT 707.5500 85.9500 709.5500 87.9500 ;
        RECT 715.7000 85.9500 717.7000 87.9500 ;
        RECT 723.8500 85.9500 725.8500 87.9500 ;
        RECT 732.0000 85.9500 734.0000 87.9500 ;
        RECT 732.0000 78.8550 734.0000 80.8550 ;
        RECT 723.8500 78.8550 725.8500 80.8550 ;
        RECT 715.7000 78.8550 717.7000 80.8550 ;
        RECT 707.5500 78.8550 709.5500 80.8550 ;
        RECT 732.0000 71.7600 734.0000 73.7600 ;
        RECT 723.8500 71.7600 725.8500 73.7600 ;
        RECT 715.7000 71.7600 717.7000 73.7600 ;
        RECT 707.5500 71.7600 709.5500 73.7600 ;
        RECT 707.5500 93.0450 709.5500 95.0450 ;
        RECT 715.7000 93.0450 717.7000 95.0450 ;
        RECT 723.8500 93.0450 725.8500 95.0450 ;
        RECT 732.0000 93.0450 734.0000 95.0450 ;
        RECT 707.5500 100.1400 709.5500 102.1400 ;
        RECT 715.7000 100.1400 717.7000 102.1400 ;
        RECT 723.8500 100.1400 725.8500 102.1400 ;
        RECT 732.0000 100.1400 734.0000 102.1400 ;
        RECT 740.1500 85.9500 742.1500 87.9500 ;
        RECT 748.3000 85.9500 750.3000 87.9500 ;
        RECT 756.4500 85.9500 758.4500 87.9500 ;
        RECT 764.6000 85.9500 766.6000 87.9500 ;
        RECT 764.6000 78.8550 766.6000 80.8550 ;
        RECT 756.4500 78.8550 758.4500 80.8550 ;
        RECT 748.3000 78.8550 750.3000 80.8550 ;
        RECT 740.1500 78.8550 742.1500 80.8550 ;
        RECT 764.6000 71.7600 766.6000 73.7600 ;
        RECT 756.4500 71.7600 758.4500 73.7600 ;
        RECT 748.3000 71.7600 750.3000 73.7600 ;
        RECT 740.1500 71.7600 742.1500 73.7600 ;
        RECT 740.1500 93.0450 742.1500 95.0450 ;
        RECT 748.3000 93.0450 750.3000 95.0450 ;
        RECT 756.4500 93.0450 758.4500 95.0450 ;
        RECT 764.6000 93.0450 766.6000 95.0450 ;
        RECT 740.1500 100.1400 742.1500 102.1400 ;
        RECT 748.3000 100.1400 750.3000 102.1400 ;
        RECT 756.4500 100.1400 758.4500 102.1400 ;
        RECT 764.6000 100.1400 766.6000 102.1400 ;
        RECT 707.5500 121.4250 709.5500 123.4250 ;
        RECT 715.7000 121.4250 717.7000 123.4250 ;
        RECT 723.8500 121.4250 725.8500 123.4250 ;
        RECT 732.0000 121.4250 734.0000 123.4250 ;
        RECT 732.0000 114.3300 734.0000 116.3300 ;
        RECT 723.8500 114.3300 725.8500 116.3300 ;
        RECT 715.7000 114.3300 717.7000 116.3300 ;
        RECT 707.5500 114.3300 709.5500 116.3300 ;
        RECT 732.0000 107.2350 734.0000 109.2350 ;
        RECT 723.8500 107.2350 725.8500 109.2350 ;
        RECT 715.7000 107.2350 717.7000 109.2350 ;
        RECT 707.5500 107.2350 709.5500 109.2350 ;
        RECT 707.5500 128.5200 709.5500 130.5200 ;
        RECT 715.7000 128.5200 717.7000 130.5200 ;
        RECT 723.8500 128.5200 725.8500 130.5200 ;
        RECT 732.0000 128.5200 734.0000 130.5200 ;
        RECT 707.5500 135.6150 709.5500 137.6150 ;
        RECT 715.7000 135.6150 717.7000 137.6150 ;
        RECT 723.8500 135.6150 725.8500 137.6150 ;
        RECT 732.0000 135.6150 734.0000 137.6150 ;
        RECT 740.1500 121.4250 742.1500 123.4250 ;
        RECT 748.3000 121.4250 750.3000 123.4250 ;
        RECT 756.4500 121.4250 758.4500 123.4250 ;
        RECT 764.6000 121.4250 766.6000 123.4250 ;
        RECT 764.6000 114.3300 766.6000 116.3300 ;
        RECT 756.4500 114.3300 758.4500 116.3300 ;
        RECT 748.3000 114.3300 750.3000 116.3300 ;
        RECT 740.1500 114.3300 742.1500 116.3300 ;
        RECT 764.6000 107.2350 766.6000 109.2350 ;
        RECT 756.4500 107.2350 758.4500 109.2350 ;
        RECT 748.3000 107.2350 750.3000 109.2350 ;
        RECT 740.1500 107.2350 742.1500 109.2350 ;
        RECT 740.1500 128.5200 742.1500 130.5200 ;
        RECT 748.3000 128.5200 750.3000 130.5200 ;
        RECT 756.4500 128.5200 758.4500 130.5200 ;
        RECT 764.6000 128.5200 766.6000 130.5200 ;
        RECT 740.1500 135.6150 742.1500 137.6150 ;
        RECT 748.3000 135.6150 750.3000 137.6150 ;
        RECT 756.4500 135.6150 758.4500 137.6150 ;
        RECT 764.6000 135.6150 766.6000 137.6150 ;
        RECT 772.7500 85.9500 774.7500 87.9500 ;
        RECT 780.9000 85.9500 782.9000 87.9500 ;
        RECT 789.0500 85.9500 791.0500 87.9500 ;
        RECT 797.2000 85.9500 799.2000 87.9500 ;
        RECT 797.2000 78.8550 799.2000 80.8550 ;
        RECT 789.0500 78.8550 791.0500 80.8550 ;
        RECT 780.9000 78.8550 782.9000 80.8550 ;
        RECT 772.7500 78.8550 774.7500 80.8550 ;
        RECT 797.2000 71.7600 799.2000 73.7600 ;
        RECT 789.0500 71.7600 791.0500 73.7600 ;
        RECT 780.9000 71.7600 782.9000 73.7600 ;
        RECT 772.7500 71.7600 774.7500 73.7600 ;
        RECT 772.7500 93.0450 774.7500 95.0450 ;
        RECT 780.9000 93.0450 782.9000 95.0450 ;
        RECT 789.0500 93.0450 791.0500 95.0450 ;
        RECT 797.2000 93.0450 799.2000 95.0450 ;
        RECT 772.7500 100.1400 774.7500 102.1400 ;
        RECT 780.9000 100.1400 782.9000 102.1400 ;
        RECT 789.0500 100.1400 791.0500 102.1400 ;
        RECT 797.2000 100.1400 799.2000 102.1400 ;
        RECT 805.3500 85.9500 807.3500 87.9500 ;
        RECT 813.5000 85.9500 815.5000 87.9500 ;
        RECT 821.6500 85.9500 823.6500 87.9500 ;
        RECT 829.8000 85.9500 831.8000 87.9500 ;
        RECT 837.9500 85.9500 839.9500 87.9500 ;
        RECT 837.9500 71.7600 839.9500 73.7600 ;
        RECT 829.8000 71.7600 831.8000 73.7600 ;
        RECT 821.6500 71.7600 823.6500 73.7600 ;
        RECT 813.5000 71.7600 815.5000 73.7600 ;
        RECT 805.3500 71.7600 807.3500 73.7600 ;
        RECT 805.3500 78.8550 807.3500 80.8550 ;
        RECT 813.5000 78.8550 815.5000 80.8550 ;
        RECT 821.6500 78.8550 823.6500 80.8550 ;
        RECT 829.8000 78.8550 831.8000 80.8550 ;
        RECT 837.9500 78.8550 839.9500 80.8550 ;
        RECT 805.3500 93.0450 807.3500 95.0450 ;
        RECT 813.5000 93.0450 815.5000 95.0450 ;
        RECT 821.6500 93.0450 823.6500 95.0450 ;
        RECT 829.8000 93.0450 831.8000 95.0450 ;
        RECT 837.9500 93.0450 839.9500 95.0450 ;
        RECT 805.3500 100.1400 807.3500 102.1400 ;
        RECT 813.5000 100.1400 815.5000 102.1400 ;
        RECT 821.6500 100.1400 823.6500 102.1400 ;
        RECT 829.8000 100.1400 831.8000 102.1400 ;
        RECT 837.9500 100.1400 839.9500 102.1400 ;
        RECT 772.7500 121.4250 774.7500 123.4250 ;
        RECT 780.9000 121.4250 782.9000 123.4250 ;
        RECT 789.0500 121.4250 791.0500 123.4250 ;
        RECT 797.2000 121.4250 799.2000 123.4250 ;
        RECT 797.2000 114.3300 799.2000 116.3300 ;
        RECT 789.0500 114.3300 791.0500 116.3300 ;
        RECT 780.9000 114.3300 782.9000 116.3300 ;
        RECT 772.7500 114.3300 774.7500 116.3300 ;
        RECT 797.2000 107.2350 799.2000 109.2350 ;
        RECT 789.0500 107.2350 791.0500 109.2350 ;
        RECT 780.9000 107.2350 782.9000 109.2350 ;
        RECT 772.7500 107.2350 774.7500 109.2350 ;
        RECT 772.7500 128.5200 774.7500 130.5200 ;
        RECT 780.9000 128.5200 782.9000 130.5200 ;
        RECT 789.0500 128.5200 791.0500 130.5200 ;
        RECT 797.2000 128.5200 799.2000 130.5200 ;
        RECT 772.7500 135.6150 774.7500 137.6150 ;
        RECT 780.9000 135.6150 782.9000 137.6150 ;
        RECT 789.0500 135.6150 791.0500 137.6150 ;
        RECT 797.2000 135.6150 799.2000 137.6150 ;
        RECT 805.3500 121.4250 807.3500 123.4250 ;
        RECT 813.5000 121.4250 815.5000 123.4250 ;
        RECT 821.6500 121.4250 823.6500 123.4250 ;
        RECT 829.8000 121.4250 831.8000 123.4250 ;
        RECT 837.9500 121.4250 839.9500 123.4250 ;
        RECT 837.9500 107.2350 839.9500 109.2350 ;
        RECT 829.8000 107.2350 831.8000 109.2350 ;
        RECT 821.6500 107.2350 823.6500 109.2350 ;
        RECT 813.5000 107.2350 815.5000 109.2350 ;
        RECT 805.3500 107.2350 807.3500 109.2350 ;
        RECT 805.3500 114.3300 807.3500 116.3300 ;
        RECT 813.5000 114.3300 815.5000 116.3300 ;
        RECT 821.6500 114.3300 823.6500 116.3300 ;
        RECT 829.8000 114.3300 831.8000 116.3300 ;
        RECT 837.9500 114.3300 839.9500 116.3300 ;
        RECT 805.3500 128.5200 807.3500 130.5200 ;
        RECT 813.5000 128.5200 815.5000 130.5200 ;
        RECT 821.6500 128.5200 823.6500 130.5200 ;
        RECT 829.8000 128.5200 831.8000 130.5200 ;
        RECT 837.9500 128.5200 839.9500 130.5200 ;
        RECT 805.3500 135.6150 807.3500 137.6150 ;
        RECT 813.5000 135.6150 815.5000 137.6150 ;
        RECT 821.6500 135.6150 823.6500 137.6150 ;
        RECT 829.8000 135.6150 831.8000 137.6150 ;
        RECT 837.9500 135.6150 839.9500 137.6150 ;
        RECT 699.4000 206.5650 701.4000 208.5650 ;
        RECT 699.4000 199.4700 701.4000 201.4700 ;
        RECT 699.4000 192.3750 701.4000 194.3750 ;
        RECT 699.4000 185.2800 701.4000 187.2800 ;
        RECT 699.4000 178.1850 701.4000 180.1850 ;
        RECT 699.4000 171.0900 701.4000 173.0900 ;
        RECT 699.4000 163.9950 701.4000 165.9950 ;
        RECT 699.4000 156.9000 701.4000 158.9000 ;
        RECT 699.4000 149.8050 701.4000 151.8050 ;
        RECT 699.4000 142.7100 701.4000 144.7100 ;
        RECT 699.4000 213.6600 701.4000 215.6600 ;
        RECT 699.4000 220.7550 701.4000 222.7550 ;
        RECT 699.4000 227.8500 701.4000 229.8500 ;
        RECT 699.4000 234.9450 701.4000 236.9450 ;
        RECT 699.4000 242.0400 701.4000 244.0400 ;
        RECT 699.4000 249.1350 701.4000 251.1350 ;
        RECT 699.4000 256.2300 701.4000 258.2300 ;
        RECT 699.4000 263.3250 701.4000 265.3250 ;
        RECT 699.4000 270.4200 701.4000 272.4200 ;
        RECT 699.4000 277.5150 701.4000 279.5150 ;
        RECT 593.4500 142.7100 595.4500 144.7100 ;
        RECT 593.4500 149.8050 595.4500 151.8050 ;
        RECT 593.4500 156.9000 595.4500 158.9000 ;
        RECT 593.4500 163.9950 595.4500 165.9950 ;
        RECT 593.4500 171.0900 595.4500 173.0900 ;
        RECT 560.8500 156.9000 562.8500 158.9000 ;
        RECT 569.0000 156.9000 571.0000 158.9000 ;
        RECT 577.1500 156.9000 579.1500 158.9000 ;
        RECT 585.3000 156.9000 587.3000 158.9000 ;
        RECT 585.3000 149.8050 587.3000 151.8050 ;
        RECT 577.1500 149.8050 579.1500 151.8050 ;
        RECT 569.0000 149.8050 571.0000 151.8050 ;
        RECT 560.8500 149.8050 562.8500 151.8050 ;
        RECT 585.3000 142.7100 587.3000 144.7100 ;
        RECT 577.1500 142.7100 579.1500 144.7100 ;
        RECT 569.0000 142.7100 571.0000 144.7100 ;
        RECT 560.8500 142.7100 562.8500 144.7100 ;
        RECT 560.8500 163.9950 562.8500 165.9950 ;
        RECT 569.0000 163.9950 571.0000 165.9950 ;
        RECT 577.1500 163.9950 579.1500 165.9950 ;
        RECT 585.3000 163.9950 587.3000 165.9950 ;
        RECT 560.8500 171.0900 562.8500 173.0900 ;
        RECT 569.0000 171.0900 571.0000 173.0900 ;
        RECT 577.1500 171.0900 579.1500 173.0900 ;
        RECT 585.3000 171.0900 587.3000 173.0900 ;
        RECT 601.6000 156.9000 603.6000 158.9000 ;
        RECT 609.7500 156.9000 611.7500 158.9000 ;
        RECT 617.9000 156.9000 619.9000 158.9000 ;
        RECT 626.0500 156.9000 628.0500 158.9000 ;
        RECT 626.0500 149.8050 628.0500 151.8050 ;
        RECT 617.9000 149.8050 619.9000 151.8050 ;
        RECT 609.7500 149.8050 611.7500 151.8050 ;
        RECT 601.6000 149.8050 603.6000 151.8050 ;
        RECT 626.0500 142.7100 628.0500 144.7100 ;
        RECT 617.9000 142.7100 619.9000 144.7100 ;
        RECT 609.7500 142.7100 611.7500 144.7100 ;
        RECT 601.6000 142.7100 603.6000 144.7100 ;
        RECT 601.6000 163.9950 603.6000 165.9950 ;
        RECT 609.7500 163.9950 611.7500 165.9950 ;
        RECT 617.9000 163.9950 619.9000 165.9950 ;
        RECT 626.0500 163.9950 628.0500 165.9950 ;
        RECT 601.6000 171.0900 603.6000 173.0900 ;
        RECT 609.7500 171.0900 611.7500 173.0900 ;
        RECT 617.9000 171.0900 619.9000 173.0900 ;
        RECT 626.0500 171.0900 628.0500 173.0900 ;
        RECT 593.4500 178.1850 595.4500 180.1850 ;
        RECT 593.4500 185.2800 595.4500 187.2800 ;
        RECT 593.4500 192.3750 595.4500 194.3750 ;
        RECT 593.4500 199.4700 595.4500 201.4700 ;
        RECT 593.4500 206.5650 595.4500 208.5650 ;
        RECT 560.8500 192.3750 562.8500 194.3750 ;
        RECT 569.0000 192.3750 571.0000 194.3750 ;
        RECT 577.1500 192.3750 579.1500 194.3750 ;
        RECT 585.3000 192.3750 587.3000 194.3750 ;
        RECT 585.3000 185.2800 587.3000 187.2800 ;
        RECT 577.1500 185.2800 579.1500 187.2800 ;
        RECT 569.0000 185.2800 571.0000 187.2800 ;
        RECT 560.8500 185.2800 562.8500 187.2800 ;
        RECT 585.3000 178.1850 587.3000 180.1850 ;
        RECT 577.1500 178.1850 579.1500 180.1850 ;
        RECT 569.0000 178.1850 571.0000 180.1850 ;
        RECT 560.8500 178.1850 562.8500 180.1850 ;
        RECT 560.8500 199.4700 562.8500 201.4700 ;
        RECT 569.0000 199.4700 571.0000 201.4700 ;
        RECT 577.1500 199.4700 579.1500 201.4700 ;
        RECT 585.3000 199.4700 587.3000 201.4700 ;
        RECT 560.8500 206.5650 562.8500 208.5650 ;
        RECT 569.0000 206.5650 571.0000 208.5650 ;
        RECT 577.1500 206.5650 579.1500 208.5650 ;
        RECT 585.3000 206.5650 587.3000 208.5650 ;
        RECT 601.6000 192.3750 603.6000 194.3750 ;
        RECT 609.7500 192.3750 611.7500 194.3750 ;
        RECT 617.9000 192.3750 619.9000 194.3750 ;
        RECT 626.0500 192.3750 628.0500 194.3750 ;
        RECT 626.0500 185.2800 628.0500 187.2800 ;
        RECT 617.9000 185.2800 619.9000 187.2800 ;
        RECT 609.7500 185.2800 611.7500 187.2800 ;
        RECT 601.6000 185.2800 603.6000 187.2800 ;
        RECT 626.0500 178.1850 628.0500 180.1850 ;
        RECT 617.9000 178.1850 619.9000 180.1850 ;
        RECT 609.7500 178.1850 611.7500 180.1850 ;
        RECT 601.6000 178.1850 603.6000 180.1850 ;
        RECT 601.6000 199.4700 603.6000 201.4700 ;
        RECT 609.7500 199.4700 611.7500 201.4700 ;
        RECT 617.9000 199.4700 619.9000 201.4700 ;
        RECT 626.0500 199.4700 628.0500 201.4700 ;
        RECT 601.6000 206.5650 603.6000 208.5650 ;
        RECT 609.7500 206.5650 611.7500 208.5650 ;
        RECT 617.9000 206.5650 619.9000 208.5650 ;
        RECT 626.0500 206.5650 628.0500 208.5650 ;
        RECT 634.2000 156.9000 636.2000 158.9000 ;
        RECT 642.3500 156.9000 644.3500 158.9000 ;
        RECT 650.5000 156.9000 652.5000 158.9000 ;
        RECT 658.6500 156.9000 660.6500 158.9000 ;
        RECT 658.6500 149.8050 660.6500 151.8050 ;
        RECT 650.5000 149.8050 652.5000 151.8050 ;
        RECT 642.3500 149.8050 644.3500 151.8050 ;
        RECT 634.2000 149.8050 636.2000 151.8050 ;
        RECT 658.6500 142.7100 660.6500 144.7100 ;
        RECT 650.5000 142.7100 652.5000 144.7100 ;
        RECT 642.3500 142.7100 644.3500 144.7100 ;
        RECT 634.2000 142.7100 636.2000 144.7100 ;
        RECT 634.2000 163.9950 636.2000 165.9950 ;
        RECT 642.3500 163.9950 644.3500 165.9950 ;
        RECT 650.5000 163.9950 652.5000 165.9950 ;
        RECT 658.6500 163.9950 660.6500 165.9950 ;
        RECT 634.2000 171.0900 636.2000 173.0900 ;
        RECT 642.3500 171.0900 644.3500 173.0900 ;
        RECT 650.5000 171.0900 652.5000 173.0900 ;
        RECT 658.6500 171.0900 660.6500 173.0900 ;
        RECT 666.8000 156.9000 668.8000 158.9000 ;
        RECT 674.9500 156.9000 676.9500 158.9000 ;
        RECT 683.1000 156.9000 685.1000 158.9000 ;
        RECT 691.2500 156.9000 693.2500 158.9000 ;
        RECT 691.2500 149.8050 693.2500 151.8050 ;
        RECT 683.1000 149.8050 685.1000 151.8050 ;
        RECT 674.9500 149.8050 676.9500 151.8050 ;
        RECT 666.8000 149.8050 668.8000 151.8050 ;
        RECT 691.2500 142.7100 693.2500 144.7100 ;
        RECT 683.1000 142.7100 685.1000 144.7100 ;
        RECT 674.9500 142.7100 676.9500 144.7100 ;
        RECT 666.8000 142.7100 668.8000 144.7100 ;
        RECT 666.8000 163.9950 668.8000 165.9950 ;
        RECT 674.9500 163.9950 676.9500 165.9950 ;
        RECT 683.1000 163.9950 685.1000 165.9950 ;
        RECT 691.2500 163.9950 693.2500 165.9950 ;
        RECT 666.8000 171.0900 668.8000 173.0900 ;
        RECT 674.9500 171.0900 676.9500 173.0900 ;
        RECT 683.1000 171.0900 685.1000 173.0900 ;
        RECT 691.2500 171.0900 693.2500 173.0900 ;
        RECT 634.2000 192.3750 636.2000 194.3750 ;
        RECT 642.3500 192.3750 644.3500 194.3750 ;
        RECT 650.5000 192.3750 652.5000 194.3750 ;
        RECT 658.6500 192.3750 660.6500 194.3750 ;
        RECT 658.6500 185.2800 660.6500 187.2800 ;
        RECT 650.5000 185.2800 652.5000 187.2800 ;
        RECT 642.3500 185.2800 644.3500 187.2800 ;
        RECT 634.2000 185.2800 636.2000 187.2800 ;
        RECT 658.6500 178.1850 660.6500 180.1850 ;
        RECT 650.5000 178.1850 652.5000 180.1850 ;
        RECT 642.3500 178.1850 644.3500 180.1850 ;
        RECT 634.2000 178.1850 636.2000 180.1850 ;
        RECT 634.2000 199.4700 636.2000 201.4700 ;
        RECT 642.3500 199.4700 644.3500 201.4700 ;
        RECT 650.5000 199.4700 652.5000 201.4700 ;
        RECT 658.6500 199.4700 660.6500 201.4700 ;
        RECT 634.2000 206.5650 636.2000 208.5650 ;
        RECT 642.3500 206.5650 644.3500 208.5650 ;
        RECT 650.5000 206.5650 652.5000 208.5650 ;
        RECT 658.6500 206.5650 660.6500 208.5650 ;
        RECT 666.8000 192.3750 668.8000 194.3750 ;
        RECT 674.9500 192.3750 676.9500 194.3750 ;
        RECT 683.1000 192.3750 685.1000 194.3750 ;
        RECT 691.2500 192.3750 693.2500 194.3750 ;
        RECT 691.2500 185.2800 693.2500 187.2800 ;
        RECT 683.1000 185.2800 685.1000 187.2800 ;
        RECT 674.9500 185.2800 676.9500 187.2800 ;
        RECT 666.8000 185.2800 668.8000 187.2800 ;
        RECT 691.2500 178.1850 693.2500 180.1850 ;
        RECT 683.1000 178.1850 685.1000 180.1850 ;
        RECT 674.9500 178.1850 676.9500 180.1850 ;
        RECT 666.8000 178.1850 668.8000 180.1850 ;
        RECT 666.8000 199.4700 668.8000 201.4700 ;
        RECT 674.9500 199.4700 676.9500 201.4700 ;
        RECT 683.1000 199.4700 685.1000 201.4700 ;
        RECT 691.2500 199.4700 693.2500 201.4700 ;
        RECT 666.8000 206.5650 668.8000 208.5650 ;
        RECT 674.9500 206.5650 676.9500 208.5650 ;
        RECT 683.1000 206.5650 685.1000 208.5650 ;
        RECT 691.2500 206.5650 693.2500 208.5650 ;
        RECT 593.4500 213.6600 595.4500 215.6600 ;
        RECT 593.4500 220.7550 595.4500 222.7550 ;
        RECT 593.4500 227.8500 595.4500 229.8500 ;
        RECT 593.4500 234.9450 595.4500 236.9450 ;
        RECT 593.4500 242.0400 595.4500 244.0400 ;
        RECT 585.3000 220.7550 587.3000 222.7550 ;
        RECT 577.1500 220.7550 579.1500 222.7550 ;
        RECT 569.0000 220.7550 571.0000 222.7550 ;
        RECT 560.8500 220.7550 562.8500 222.7550 ;
        RECT 585.3000 213.6600 587.3000 215.6600 ;
        RECT 577.1500 213.6600 579.1500 215.6600 ;
        RECT 569.0000 213.6600 571.0000 215.6600 ;
        RECT 560.8500 213.6600 562.8500 215.6600 ;
        RECT 569.0000 227.8500 571.0000 229.8500 ;
        RECT 560.8500 227.8500 562.8500 229.8500 ;
        RECT 577.1500 227.8500 579.1500 229.8500 ;
        RECT 585.3000 227.8500 587.3000 229.8500 ;
        RECT 560.8500 234.9450 562.8500 236.9450 ;
        RECT 569.0000 234.9450 571.0000 236.9450 ;
        RECT 577.1500 234.9450 579.1500 236.9450 ;
        RECT 585.3000 234.9450 587.3000 236.9450 ;
        RECT 560.8500 242.0400 562.8500 244.0400 ;
        RECT 569.0000 242.0400 571.0000 244.0400 ;
        RECT 577.1500 242.0400 579.1500 244.0400 ;
        RECT 585.3000 242.0400 587.3000 244.0400 ;
        RECT 626.0500 220.7550 628.0500 222.7550 ;
        RECT 617.9000 220.7550 619.9000 222.7550 ;
        RECT 609.7500 220.7550 611.7500 222.7550 ;
        RECT 601.6000 220.7550 603.6000 222.7550 ;
        RECT 626.0500 213.6600 628.0500 215.6600 ;
        RECT 617.9000 213.6600 619.9000 215.6600 ;
        RECT 609.7500 213.6600 611.7500 215.6600 ;
        RECT 601.6000 213.6600 603.6000 215.6600 ;
        RECT 609.7500 227.8500 611.7500 229.8500 ;
        RECT 601.6000 227.8500 603.6000 229.8500 ;
        RECT 617.9000 227.8500 619.9000 229.8500 ;
        RECT 626.0500 227.8500 628.0500 229.8500 ;
        RECT 601.6000 234.9450 603.6000 236.9450 ;
        RECT 609.7500 234.9450 611.7500 236.9450 ;
        RECT 617.9000 234.9450 619.9000 236.9450 ;
        RECT 626.0500 234.9450 628.0500 236.9450 ;
        RECT 601.6000 242.0400 603.6000 244.0400 ;
        RECT 609.7500 242.0400 611.7500 244.0400 ;
        RECT 617.9000 242.0400 619.9000 244.0400 ;
        RECT 626.0500 242.0400 628.0500 244.0400 ;
        RECT 593.4500 249.1350 595.4500 251.1350 ;
        RECT 593.4500 256.2300 595.4500 258.2300 ;
        RECT 593.4500 263.3250 595.4500 265.3250 ;
        RECT 593.4500 270.4200 595.4500 272.4200 ;
        RECT 593.4500 277.5150 595.4500 279.5150 ;
        RECT 585.3000 256.2300 587.3000 258.2300 ;
        RECT 577.1500 256.2300 579.1500 258.2300 ;
        RECT 569.0000 256.2300 571.0000 258.2300 ;
        RECT 560.8500 256.2300 562.8500 258.2300 ;
        RECT 585.3000 249.1350 587.3000 251.1350 ;
        RECT 577.1500 249.1350 579.1500 251.1350 ;
        RECT 569.0000 249.1350 571.0000 251.1350 ;
        RECT 560.8500 249.1350 562.8500 251.1350 ;
        RECT 569.0000 263.3250 571.0000 265.3250 ;
        RECT 560.8500 263.3250 562.8500 265.3250 ;
        RECT 577.1500 263.3250 579.1500 265.3250 ;
        RECT 585.3000 263.3250 587.3000 265.3250 ;
        RECT 560.8500 270.4200 562.8500 272.4200 ;
        RECT 569.0000 270.4200 571.0000 272.4200 ;
        RECT 577.1500 270.4200 579.1500 272.4200 ;
        RECT 585.3000 270.4200 587.3000 272.4200 ;
        RECT 560.8500 277.5150 562.8500 279.5150 ;
        RECT 569.0000 277.5150 571.0000 279.5150 ;
        RECT 577.1500 277.5150 579.1500 279.5150 ;
        RECT 585.3000 277.5150 587.3000 279.5150 ;
        RECT 626.0500 256.2300 628.0500 258.2300 ;
        RECT 617.9000 256.2300 619.9000 258.2300 ;
        RECT 609.7500 256.2300 611.7500 258.2300 ;
        RECT 601.6000 256.2300 603.6000 258.2300 ;
        RECT 626.0500 249.1350 628.0500 251.1350 ;
        RECT 617.9000 249.1350 619.9000 251.1350 ;
        RECT 609.7500 249.1350 611.7500 251.1350 ;
        RECT 601.6000 249.1350 603.6000 251.1350 ;
        RECT 609.7500 263.3250 611.7500 265.3250 ;
        RECT 601.6000 263.3250 603.6000 265.3250 ;
        RECT 617.9000 263.3250 619.9000 265.3250 ;
        RECT 626.0500 263.3250 628.0500 265.3250 ;
        RECT 601.6000 270.4200 603.6000 272.4200 ;
        RECT 609.7500 270.4200 611.7500 272.4200 ;
        RECT 617.9000 270.4200 619.9000 272.4200 ;
        RECT 626.0500 270.4200 628.0500 272.4200 ;
        RECT 601.6000 277.5150 603.6000 279.5150 ;
        RECT 609.7500 277.5150 611.7500 279.5150 ;
        RECT 617.9000 277.5150 619.9000 279.5150 ;
        RECT 626.0500 277.5150 628.0500 279.5150 ;
        RECT 658.6500 220.7550 660.6500 222.7550 ;
        RECT 650.5000 220.7550 652.5000 222.7550 ;
        RECT 642.3500 220.7550 644.3500 222.7550 ;
        RECT 634.2000 220.7550 636.2000 222.7550 ;
        RECT 658.6500 213.6600 660.6500 215.6600 ;
        RECT 650.5000 213.6600 652.5000 215.6600 ;
        RECT 642.3500 213.6600 644.3500 215.6600 ;
        RECT 634.2000 213.6600 636.2000 215.6600 ;
        RECT 642.3500 227.8500 644.3500 229.8500 ;
        RECT 634.2000 227.8500 636.2000 229.8500 ;
        RECT 650.5000 227.8500 652.5000 229.8500 ;
        RECT 658.6500 227.8500 660.6500 229.8500 ;
        RECT 634.2000 234.9450 636.2000 236.9450 ;
        RECT 642.3500 234.9450 644.3500 236.9450 ;
        RECT 650.5000 234.9450 652.5000 236.9450 ;
        RECT 658.6500 234.9450 660.6500 236.9450 ;
        RECT 634.2000 242.0400 636.2000 244.0400 ;
        RECT 642.3500 242.0400 644.3500 244.0400 ;
        RECT 650.5000 242.0400 652.5000 244.0400 ;
        RECT 658.6500 242.0400 660.6500 244.0400 ;
        RECT 691.2500 220.7550 693.2500 222.7550 ;
        RECT 683.1000 220.7550 685.1000 222.7550 ;
        RECT 674.9500 220.7550 676.9500 222.7550 ;
        RECT 666.8000 220.7550 668.8000 222.7550 ;
        RECT 691.2500 213.6600 693.2500 215.6600 ;
        RECT 683.1000 213.6600 685.1000 215.6600 ;
        RECT 674.9500 213.6600 676.9500 215.6600 ;
        RECT 666.8000 213.6600 668.8000 215.6600 ;
        RECT 674.9500 227.8500 676.9500 229.8500 ;
        RECT 666.8000 227.8500 668.8000 229.8500 ;
        RECT 683.1000 227.8500 685.1000 229.8500 ;
        RECT 691.2500 227.8500 693.2500 229.8500 ;
        RECT 666.8000 234.9450 668.8000 236.9450 ;
        RECT 674.9500 234.9450 676.9500 236.9450 ;
        RECT 683.1000 234.9450 685.1000 236.9450 ;
        RECT 691.2500 234.9450 693.2500 236.9450 ;
        RECT 666.8000 242.0400 668.8000 244.0400 ;
        RECT 674.9500 242.0400 676.9500 244.0400 ;
        RECT 683.1000 242.0400 685.1000 244.0400 ;
        RECT 691.2500 242.0400 693.2500 244.0400 ;
        RECT 658.6500 256.2300 660.6500 258.2300 ;
        RECT 650.5000 256.2300 652.5000 258.2300 ;
        RECT 642.3500 256.2300 644.3500 258.2300 ;
        RECT 634.2000 256.2300 636.2000 258.2300 ;
        RECT 658.6500 249.1350 660.6500 251.1350 ;
        RECT 650.5000 249.1350 652.5000 251.1350 ;
        RECT 642.3500 249.1350 644.3500 251.1350 ;
        RECT 634.2000 249.1350 636.2000 251.1350 ;
        RECT 642.3500 263.3250 644.3500 265.3250 ;
        RECT 634.2000 263.3250 636.2000 265.3250 ;
        RECT 650.5000 263.3250 652.5000 265.3250 ;
        RECT 658.6500 263.3250 660.6500 265.3250 ;
        RECT 634.2000 270.4200 636.2000 272.4200 ;
        RECT 642.3500 270.4200 644.3500 272.4200 ;
        RECT 650.5000 270.4200 652.5000 272.4200 ;
        RECT 658.6500 270.4200 660.6500 272.4200 ;
        RECT 634.2000 277.5150 636.2000 279.5150 ;
        RECT 642.3500 277.5150 644.3500 279.5150 ;
        RECT 650.5000 277.5150 652.5000 279.5150 ;
        RECT 658.6500 277.5150 660.6500 279.5150 ;
        RECT 691.2500 256.2300 693.2500 258.2300 ;
        RECT 683.1000 256.2300 685.1000 258.2300 ;
        RECT 674.9500 256.2300 676.9500 258.2300 ;
        RECT 666.8000 256.2300 668.8000 258.2300 ;
        RECT 691.2500 249.1350 693.2500 251.1350 ;
        RECT 683.1000 249.1350 685.1000 251.1350 ;
        RECT 674.9500 249.1350 676.9500 251.1350 ;
        RECT 666.8000 249.1350 668.8000 251.1350 ;
        RECT 674.9500 263.3250 676.9500 265.3250 ;
        RECT 666.8000 263.3250 668.8000 265.3250 ;
        RECT 683.1000 263.3250 685.1000 265.3250 ;
        RECT 691.2500 263.3250 693.2500 265.3250 ;
        RECT 666.8000 270.4200 668.8000 272.4200 ;
        RECT 674.9500 270.4200 676.9500 272.4200 ;
        RECT 683.1000 270.4200 685.1000 272.4200 ;
        RECT 691.2500 270.4200 693.2500 272.4200 ;
        RECT 666.8000 277.5150 668.8000 279.5150 ;
        RECT 674.9500 277.5150 676.9500 279.5150 ;
        RECT 683.1000 277.5150 685.1000 279.5150 ;
        RECT 691.2500 277.5150 693.2500 279.5150 ;
        RECT 707.5500 156.9000 709.5500 158.9000 ;
        RECT 715.7000 156.9000 717.7000 158.9000 ;
        RECT 723.8500 156.9000 725.8500 158.9000 ;
        RECT 732.0000 156.9000 734.0000 158.9000 ;
        RECT 732.0000 149.8050 734.0000 151.8050 ;
        RECT 723.8500 149.8050 725.8500 151.8050 ;
        RECT 715.7000 149.8050 717.7000 151.8050 ;
        RECT 707.5500 149.8050 709.5500 151.8050 ;
        RECT 732.0000 142.7100 734.0000 144.7100 ;
        RECT 723.8500 142.7100 725.8500 144.7100 ;
        RECT 715.7000 142.7100 717.7000 144.7100 ;
        RECT 707.5500 142.7100 709.5500 144.7100 ;
        RECT 707.5500 163.9950 709.5500 165.9950 ;
        RECT 715.7000 163.9950 717.7000 165.9950 ;
        RECT 723.8500 163.9950 725.8500 165.9950 ;
        RECT 732.0000 163.9950 734.0000 165.9950 ;
        RECT 707.5500 171.0900 709.5500 173.0900 ;
        RECT 715.7000 171.0900 717.7000 173.0900 ;
        RECT 723.8500 171.0900 725.8500 173.0900 ;
        RECT 732.0000 171.0900 734.0000 173.0900 ;
        RECT 740.1500 156.9000 742.1500 158.9000 ;
        RECT 748.3000 156.9000 750.3000 158.9000 ;
        RECT 756.4500 156.9000 758.4500 158.9000 ;
        RECT 764.6000 156.9000 766.6000 158.9000 ;
        RECT 764.6000 149.8050 766.6000 151.8050 ;
        RECT 756.4500 149.8050 758.4500 151.8050 ;
        RECT 748.3000 149.8050 750.3000 151.8050 ;
        RECT 740.1500 149.8050 742.1500 151.8050 ;
        RECT 764.6000 142.7100 766.6000 144.7100 ;
        RECT 756.4500 142.7100 758.4500 144.7100 ;
        RECT 748.3000 142.7100 750.3000 144.7100 ;
        RECT 740.1500 142.7100 742.1500 144.7100 ;
        RECT 740.1500 163.9950 742.1500 165.9950 ;
        RECT 748.3000 163.9950 750.3000 165.9950 ;
        RECT 756.4500 163.9950 758.4500 165.9950 ;
        RECT 764.6000 163.9950 766.6000 165.9950 ;
        RECT 740.1500 171.0900 742.1500 173.0900 ;
        RECT 748.3000 171.0900 750.3000 173.0900 ;
        RECT 756.4500 171.0900 758.4500 173.0900 ;
        RECT 764.6000 171.0900 766.6000 173.0900 ;
        RECT 707.5500 192.3750 709.5500 194.3750 ;
        RECT 715.7000 192.3750 717.7000 194.3750 ;
        RECT 723.8500 192.3750 725.8500 194.3750 ;
        RECT 732.0000 192.3750 734.0000 194.3750 ;
        RECT 732.0000 185.2800 734.0000 187.2800 ;
        RECT 723.8500 185.2800 725.8500 187.2800 ;
        RECT 715.7000 185.2800 717.7000 187.2800 ;
        RECT 707.5500 185.2800 709.5500 187.2800 ;
        RECT 732.0000 178.1850 734.0000 180.1850 ;
        RECT 723.8500 178.1850 725.8500 180.1850 ;
        RECT 715.7000 178.1850 717.7000 180.1850 ;
        RECT 707.5500 178.1850 709.5500 180.1850 ;
        RECT 707.5500 199.4700 709.5500 201.4700 ;
        RECT 715.7000 199.4700 717.7000 201.4700 ;
        RECT 723.8500 199.4700 725.8500 201.4700 ;
        RECT 732.0000 199.4700 734.0000 201.4700 ;
        RECT 707.5500 206.5650 709.5500 208.5650 ;
        RECT 715.7000 206.5650 717.7000 208.5650 ;
        RECT 723.8500 206.5650 725.8500 208.5650 ;
        RECT 732.0000 206.5650 734.0000 208.5650 ;
        RECT 740.1500 192.3750 742.1500 194.3750 ;
        RECT 748.3000 192.3750 750.3000 194.3750 ;
        RECT 756.4500 192.3750 758.4500 194.3750 ;
        RECT 764.6000 192.3750 766.6000 194.3750 ;
        RECT 764.6000 185.2800 766.6000 187.2800 ;
        RECT 756.4500 185.2800 758.4500 187.2800 ;
        RECT 748.3000 185.2800 750.3000 187.2800 ;
        RECT 740.1500 185.2800 742.1500 187.2800 ;
        RECT 764.6000 178.1850 766.6000 180.1850 ;
        RECT 756.4500 178.1850 758.4500 180.1850 ;
        RECT 748.3000 178.1850 750.3000 180.1850 ;
        RECT 740.1500 178.1850 742.1500 180.1850 ;
        RECT 740.1500 199.4700 742.1500 201.4700 ;
        RECT 748.3000 199.4700 750.3000 201.4700 ;
        RECT 756.4500 199.4700 758.4500 201.4700 ;
        RECT 764.6000 199.4700 766.6000 201.4700 ;
        RECT 740.1500 206.5650 742.1500 208.5650 ;
        RECT 748.3000 206.5650 750.3000 208.5650 ;
        RECT 756.4500 206.5650 758.4500 208.5650 ;
        RECT 764.6000 206.5650 766.6000 208.5650 ;
        RECT 772.7500 156.9000 774.7500 158.9000 ;
        RECT 780.9000 156.9000 782.9000 158.9000 ;
        RECT 789.0500 156.9000 791.0500 158.9000 ;
        RECT 797.2000 156.9000 799.2000 158.9000 ;
        RECT 797.2000 149.8050 799.2000 151.8050 ;
        RECT 789.0500 149.8050 791.0500 151.8050 ;
        RECT 780.9000 149.8050 782.9000 151.8050 ;
        RECT 772.7500 149.8050 774.7500 151.8050 ;
        RECT 797.2000 142.7100 799.2000 144.7100 ;
        RECT 789.0500 142.7100 791.0500 144.7100 ;
        RECT 780.9000 142.7100 782.9000 144.7100 ;
        RECT 772.7500 142.7100 774.7500 144.7100 ;
        RECT 772.7500 163.9950 774.7500 165.9950 ;
        RECT 780.9000 163.9950 782.9000 165.9950 ;
        RECT 789.0500 163.9950 791.0500 165.9950 ;
        RECT 797.2000 163.9950 799.2000 165.9950 ;
        RECT 772.7500 171.0900 774.7500 173.0900 ;
        RECT 780.9000 171.0900 782.9000 173.0900 ;
        RECT 789.0500 171.0900 791.0500 173.0900 ;
        RECT 797.2000 171.0900 799.2000 173.0900 ;
        RECT 805.3500 156.9000 807.3500 158.9000 ;
        RECT 813.5000 156.9000 815.5000 158.9000 ;
        RECT 821.6500 156.9000 823.6500 158.9000 ;
        RECT 829.8000 156.9000 831.8000 158.9000 ;
        RECT 837.9500 156.9000 839.9500 158.9000 ;
        RECT 837.9500 142.7100 839.9500 144.7100 ;
        RECT 829.8000 142.7100 831.8000 144.7100 ;
        RECT 821.6500 142.7100 823.6500 144.7100 ;
        RECT 813.5000 142.7100 815.5000 144.7100 ;
        RECT 805.3500 142.7100 807.3500 144.7100 ;
        RECT 805.3500 149.8050 807.3500 151.8050 ;
        RECT 813.5000 149.8050 815.5000 151.8050 ;
        RECT 821.6500 149.8050 823.6500 151.8050 ;
        RECT 829.8000 149.8050 831.8000 151.8050 ;
        RECT 837.9500 149.8050 839.9500 151.8050 ;
        RECT 805.3500 163.9950 807.3500 165.9950 ;
        RECT 813.5000 163.9950 815.5000 165.9950 ;
        RECT 821.6500 163.9950 823.6500 165.9950 ;
        RECT 829.8000 163.9950 831.8000 165.9950 ;
        RECT 837.9500 163.9950 839.9500 165.9950 ;
        RECT 805.3500 171.0900 807.3500 173.0900 ;
        RECT 813.5000 171.0900 815.5000 173.0900 ;
        RECT 821.6500 171.0900 823.6500 173.0900 ;
        RECT 829.8000 171.0900 831.8000 173.0900 ;
        RECT 837.9500 171.0900 839.9500 173.0900 ;
        RECT 772.7500 192.3750 774.7500 194.3750 ;
        RECT 780.9000 192.3750 782.9000 194.3750 ;
        RECT 789.0500 192.3750 791.0500 194.3750 ;
        RECT 797.2000 192.3750 799.2000 194.3750 ;
        RECT 797.2000 185.2800 799.2000 187.2800 ;
        RECT 789.0500 185.2800 791.0500 187.2800 ;
        RECT 780.9000 185.2800 782.9000 187.2800 ;
        RECT 772.7500 185.2800 774.7500 187.2800 ;
        RECT 797.2000 178.1850 799.2000 180.1850 ;
        RECT 789.0500 178.1850 791.0500 180.1850 ;
        RECT 780.9000 178.1850 782.9000 180.1850 ;
        RECT 772.7500 178.1850 774.7500 180.1850 ;
        RECT 772.7500 199.4700 774.7500 201.4700 ;
        RECT 780.9000 199.4700 782.9000 201.4700 ;
        RECT 789.0500 199.4700 791.0500 201.4700 ;
        RECT 797.2000 199.4700 799.2000 201.4700 ;
        RECT 772.7500 206.5650 774.7500 208.5650 ;
        RECT 780.9000 206.5650 782.9000 208.5650 ;
        RECT 789.0500 206.5650 791.0500 208.5650 ;
        RECT 797.2000 206.5650 799.2000 208.5650 ;
        RECT 805.3500 192.3750 807.3500 194.3750 ;
        RECT 813.5000 192.3750 815.5000 194.3750 ;
        RECT 821.6500 192.3750 823.6500 194.3750 ;
        RECT 829.8000 192.3750 831.8000 194.3750 ;
        RECT 837.9500 192.3750 839.9500 194.3750 ;
        RECT 837.9500 178.1850 839.9500 180.1850 ;
        RECT 829.8000 178.1850 831.8000 180.1850 ;
        RECT 821.6500 178.1850 823.6500 180.1850 ;
        RECT 813.5000 178.1850 815.5000 180.1850 ;
        RECT 805.3500 178.1850 807.3500 180.1850 ;
        RECT 805.3500 185.2800 807.3500 187.2800 ;
        RECT 813.5000 185.2800 815.5000 187.2800 ;
        RECT 821.6500 185.2800 823.6500 187.2800 ;
        RECT 829.8000 185.2800 831.8000 187.2800 ;
        RECT 837.9500 185.2800 839.9500 187.2800 ;
        RECT 805.3500 199.4700 807.3500 201.4700 ;
        RECT 813.5000 199.4700 815.5000 201.4700 ;
        RECT 821.6500 199.4700 823.6500 201.4700 ;
        RECT 829.8000 199.4700 831.8000 201.4700 ;
        RECT 837.9500 199.4700 839.9500 201.4700 ;
        RECT 805.3500 206.5650 807.3500 208.5650 ;
        RECT 813.5000 206.5650 815.5000 208.5650 ;
        RECT 821.6500 206.5650 823.6500 208.5650 ;
        RECT 829.8000 206.5650 831.8000 208.5650 ;
        RECT 837.9500 206.5650 839.9500 208.5650 ;
        RECT 732.0000 220.7550 734.0000 222.7550 ;
        RECT 723.8500 220.7550 725.8500 222.7550 ;
        RECT 715.7000 220.7550 717.7000 222.7550 ;
        RECT 707.5500 220.7550 709.5500 222.7550 ;
        RECT 732.0000 213.6600 734.0000 215.6600 ;
        RECT 723.8500 213.6600 725.8500 215.6600 ;
        RECT 715.7000 213.6600 717.7000 215.6600 ;
        RECT 707.5500 213.6600 709.5500 215.6600 ;
        RECT 715.7000 227.8500 717.7000 229.8500 ;
        RECT 707.5500 227.8500 709.5500 229.8500 ;
        RECT 723.8500 227.8500 725.8500 229.8500 ;
        RECT 732.0000 227.8500 734.0000 229.8500 ;
        RECT 707.5500 234.9450 709.5500 236.9450 ;
        RECT 715.7000 234.9450 717.7000 236.9450 ;
        RECT 723.8500 234.9450 725.8500 236.9450 ;
        RECT 732.0000 234.9450 734.0000 236.9450 ;
        RECT 707.5500 242.0400 709.5500 244.0400 ;
        RECT 715.7000 242.0400 717.7000 244.0400 ;
        RECT 723.8500 242.0400 725.8500 244.0400 ;
        RECT 732.0000 242.0400 734.0000 244.0400 ;
        RECT 764.6000 220.7550 766.6000 222.7550 ;
        RECT 756.4500 220.7550 758.4500 222.7550 ;
        RECT 748.3000 220.7550 750.3000 222.7550 ;
        RECT 740.1500 220.7550 742.1500 222.7550 ;
        RECT 764.6000 213.6600 766.6000 215.6600 ;
        RECT 756.4500 213.6600 758.4500 215.6600 ;
        RECT 748.3000 213.6600 750.3000 215.6600 ;
        RECT 740.1500 213.6600 742.1500 215.6600 ;
        RECT 748.3000 227.8500 750.3000 229.8500 ;
        RECT 740.1500 227.8500 742.1500 229.8500 ;
        RECT 756.4500 227.8500 758.4500 229.8500 ;
        RECT 764.6000 227.8500 766.6000 229.8500 ;
        RECT 740.1500 234.9450 742.1500 236.9450 ;
        RECT 748.3000 234.9450 750.3000 236.9450 ;
        RECT 756.4500 234.9450 758.4500 236.9450 ;
        RECT 764.6000 234.9450 766.6000 236.9450 ;
        RECT 740.1500 242.0400 742.1500 244.0400 ;
        RECT 748.3000 242.0400 750.3000 244.0400 ;
        RECT 756.4500 242.0400 758.4500 244.0400 ;
        RECT 764.6000 242.0400 766.6000 244.0400 ;
        RECT 732.0000 256.2300 734.0000 258.2300 ;
        RECT 723.8500 256.2300 725.8500 258.2300 ;
        RECT 715.7000 256.2300 717.7000 258.2300 ;
        RECT 707.5500 256.2300 709.5500 258.2300 ;
        RECT 732.0000 249.1350 734.0000 251.1350 ;
        RECT 723.8500 249.1350 725.8500 251.1350 ;
        RECT 715.7000 249.1350 717.7000 251.1350 ;
        RECT 707.5500 249.1350 709.5500 251.1350 ;
        RECT 715.7000 263.3250 717.7000 265.3250 ;
        RECT 707.5500 263.3250 709.5500 265.3250 ;
        RECT 723.8500 263.3250 725.8500 265.3250 ;
        RECT 732.0000 263.3250 734.0000 265.3250 ;
        RECT 707.5500 270.4200 709.5500 272.4200 ;
        RECT 715.7000 270.4200 717.7000 272.4200 ;
        RECT 723.8500 270.4200 725.8500 272.4200 ;
        RECT 732.0000 270.4200 734.0000 272.4200 ;
        RECT 707.5500 277.5150 709.5500 279.5150 ;
        RECT 715.7000 277.5150 717.7000 279.5150 ;
        RECT 723.8500 277.5150 725.8500 279.5150 ;
        RECT 732.0000 277.5150 734.0000 279.5150 ;
        RECT 764.6000 256.2300 766.6000 258.2300 ;
        RECT 756.4500 256.2300 758.4500 258.2300 ;
        RECT 748.3000 256.2300 750.3000 258.2300 ;
        RECT 740.1500 256.2300 742.1500 258.2300 ;
        RECT 764.6000 249.1350 766.6000 251.1350 ;
        RECT 756.4500 249.1350 758.4500 251.1350 ;
        RECT 748.3000 249.1350 750.3000 251.1350 ;
        RECT 740.1500 249.1350 742.1500 251.1350 ;
        RECT 748.3000 263.3250 750.3000 265.3250 ;
        RECT 740.1500 263.3250 742.1500 265.3250 ;
        RECT 756.4500 263.3250 758.4500 265.3250 ;
        RECT 764.6000 263.3250 766.6000 265.3250 ;
        RECT 740.1500 270.4200 742.1500 272.4200 ;
        RECT 748.3000 270.4200 750.3000 272.4200 ;
        RECT 756.4500 270.4200 758.4500 272.4200 ;
        RECT 764.6000 270.4200 766.6000 272.4200 ;
        RECT 740.1500 277.5150 742.1500 279.5150 ;
        RECT 748.3000 277.5150 750.3000 279.5150 ;
        RECT 756.4500 277.5150 758.4500 279.5150 ;
        RECT 764.6000 277.5150 766.6000 279.5150 ;
        RECT 797.2000 220.7550 799.2000 222.7550 ;
        RECT 789.0500 220.7550 791.0500 222.7550 ;
        RECT 780.9000 220.7550 782.9000 222.7550 ;
        RECT 772.7500 220.7550 774.7500 222.7550 ;
        RECT 797.2000 213.6600 799.2000 215.6600 ;
        RECT 789.0500 213.6600 791.0500 215.6600 ;
        RECT 780.9000 213.6600 782.9000 215.6600 ;
        RECT 772.7500 213.6600 774.7500 215.6600 ;
        RECT 780.9000 227.8500 782.9000 229.8500 ;
        RECT 772.7500 227.8500 774.7500 229.8500 ;
        RECT 789.0500 227.8500 791.0500 229.8500 ;
        RECT 797.2000 227.8500 799.2000 229.8500 ;
        RECT 772.7500 234.9450 774.7500 236.9450 ;
        RECT 780.9000 234.9450 782.9000 236.9450 ;
        RECT 789.0500 234.9450 791.0500 236.9450 ;
        RECT 797.2000 234.9450 799.2000 236.9450 ;
        RECT 772.7500 242.0400 774.7500 244.0400 ;
        RECT 780.9000 242.0400 782.9000 244.0400 ;
        RECT 789.0500 242.0400 791.0500 244.0400 ;
        RECT 797.2000 242.0400 799.2000 244.0400 ;
        RECT 837.9500 213.6600 839.9500 215.6600 ;
        RECT 829.8000 213.6600 831.8000 215.6600 ;
        RECT 821.6500 213.6600 823.6500 215.6600 ;
        RECT 813.5000 213.6600 815.5000 215.6600 ;
        RECT 805.3500 213.6600 807.3500 215.6600 ;
        RECT 805.3500 220.7550 807.3500 222.7550 ;
        RECT 813.5000 220.7550 815.5000 222.7550 ;
        RECT 821.6500 220.7550 823.6500 222.7550 ;
        RECT 829.8000 220.7550 831.8000 222.7550 ;
        RECT 837.9500 220.7550 839.9500 222.7550 ;
        RECT 821.6500 227.8500 823.6500 229.8500 ;
        RECT 821.6500 234.9450 823.6500 236.9450 ;
        RECT 821.6500 242.0400 823.6500 244.0400 ;
        RECT 813.5000 242.0400 815.5000 244.0400 ;
        RECT 805.3500 242.0400 807.3500 244.0400 ;
        RECT 813.5000 234.9450 815.5000 236.9450 ;
        RECT 805.3500 234.9450 807.3500 236.9450 ;
        RECT 813.5000 227.8500 815.5000 229.8500 ;
        RECT 805.3500 227.8500 807.3500 229.8500 ;
        RECT 837.9500 242.0400 839.9500 244.0400 ;
        RECT 829.8000 242.0400 831.8000 244.0400 ;
        RECT 837.9500 234.9450 839.9500 236.9450 ;
        RECT 829.8000 234.9450 831.8000 236.9450 ;
        RECT 837.9500 227.8500 839.9500 229.8500 ;
        RECT 829.8000 227.8500 831.8000 229.8500 ;
        RECT 797.2000 256.2300 799.2000 258.2300 ;
        RECT 789.0500 256.2300 791.0500 258.2300 ;
        RECT 780.9000 256.2300 782.9000 258.2300 ;
        RECT 772.7500 256.2300 774.7500 258.2300 ;
        RECT 797.2000 249.1350 799.2000 251.1350 ;
        RECT 789.0500 249.1350 791.0500 251.1350 ;
        RECT 780.9000 249.1350 782.9000 251.1350 ;
        RECT 772.7500 249.1350 774.7500 251.1350 ;
        RECT 780.9000 263.3250 782.9000 265.3250 ;
        RECT 772.7500 263.3250 774.7500 265.3250 ;
        RECT 789.0500 263.3250 791.0500 265.3250 ;
        RECT 797.2000 263.3250 799.2000 265.3250 ;
        RECT 772.7500 270.4200 774.7500 272.4200 ;
        RECT 780.9000 270.4200 782.9000 272.4200 ;
        RECT 789.0500 270.4200 791.0500 272.4200 ;
        RECT 797.2000 270.4200 799.2000 272.4200 ;
        RECT 772.7500 277.5150 774.7500 279.5150 ;
        RECT 780.9000 277.5150 782.9000 279.5150 ;
        RECT 789.0500 277.5150 791.0500 279.5150 ;
        RECT 797.2000 277.5150 799.2000 279.5150 ;
        RECT 837.9500 249.1350 839.9500 251.1350 ;
        RECT 829.8000 249.1350 831.8000 251.1350 ;
        RECT 821.6500 249.1350 823.6500 251.1350 ;
        RECT 813.5000 249.1350 815.5000 251.1350 ;
        RECT 805.3500 249.1350 807.3500 251.1350 ;
        RECT 805.3500 256.2300 807.3500 258.2300 ;
        RECT 813.5000 256.2300 815.5000 258.2300 ;
        RECT 821.6500 256.2300 823.6500 258.2300 ;
        RECT 829.8000 256.2300 831.8000 258.2300 ;
        RECT 837.9500 256.2300 839.9500 258.2300 ;
        RECT 821.6500 263.3250 823.6500 265.3250 ;
        RECT 821.6500 270.4200 823.6500 272.4200 ;
        RECT 821.6500 277.5150 823.6500 279.5150 ;
        RECT 813.5000 277.5150 815.5000 279.5150 ;
        RECT 805.3500 277.5150 807.3500 279.5150 ;
        RECT 813.5000 270.4200 815.5000 272.4200 ;
        RECT 805.3500 270.4200 807.3500 272.4200 ;
        RECT 813.5000 263.3250 815.5000 265.3250 ;
        RECT 805.3500 263.3250 807.3500 265.3250 ;
        RECT 837.9500 277.5150 839.9500 279.5150 ;
        RECT 829.8000 277.5150 831.8000 279.5150 ;
        RECT 837.9500 270.4200 839.9500 272.4200 ;
        RECT 829.8000 270.4200 831.8000 272.4200 ;
        RECT 837.9500 263.3250 839.9500 265.3250 ;
        RECT 829.8000 263.3250 831.8000 265.3250 ;
        RECT 903.1500 64.6650 905.1500 66.6650 ;
        RECT 895.0000 64.6650 897.0000 66.6650 ;
        RECT 886.8500 64.6650 888.8500 66.6650 ;
        RECT 878.7000 64.6650 880.7000 66.6650 ;
        RECT 870.5500 64.6650 872.5500 66.6650 ;
        RECT 862.4000 64.6650 864.4000 66.6650 ;
        RECT 854.2500 64.6650 856.2500 66.6650 ;
        RECT 846.1000 64.6650 848.1000 66.6650 ;
        RECT 943.9000 64.6650 945.9000 66.6650 ;
        RECT 935.7500 64.6650 937.7500 66.6650 ;
        RECT 927.6000 64.6650 929.6000 66.6650 ;
        RECT 919.4500 64.6650 921.4500 66.6650 ;
        RECT 911.3000 64.6650 913.3000 66.6650 ;
        RECT 952.0500 64.6650 954.0500 66.6650 ;
        RECT 960.2000 64.6650 962.2000 66.6650 ;
        RECT 968.3500 64.6650 970.3500 66.6650 ;
        RECT 976.5000 64.6650 978.5000 66.6650 ;
        RECT 846.1000 85.9500 848.1000 87.9500 ;
        RECT 854.2500 85.9500 856.2500 87.9500 ;
        RECT 862.4000 85.9500 864.4000 87.9500 ;
        RECT 870.5500 85.9500 872.5500 87.9500 ;
        RECT 870.5500 78.8550 872.5500 80.8550 ;
        RECT 862.4000 78.8550 864.4000 80.8550 ;
        RECT 854.2500 78.8550 856.2500 80.8550 ;
        RECT 846.1000 78.8550 848.1000 80.8550 ;
        RECT 870.5500 71.7600 872.5500 73.7600 ;
        RECT 862.4000 71.7600 864.4000 73.7600 ;
        RECT 854.2500 71.7600 856.2500 73.7600 ;
        RECT 846.1000 71.7600 848.1000 73.7600 ;
        RECT 846.1000 93.0450 848.1000 95.0450 ;
        RECT 854.2500 93.0450 856.2500 95.0450 ;
        RECT 862.4000 93.0450 864.4000 95.0450 ;
        RECT 870.5500 93.0450 872.5500 95.0450 ;
        RECT 846.1000 100.1400 848.1000 102.1400 ;
        RECT 854.2500 100.1400 856.2500 102.1400 ;
        RECT 862.4000 100.1400 864.4000 102.1400 ;
        RECT 870.5500 100.1400 872.5500 102.1400 ;
        RECT 878.7000 85.9500 880.7000 87.9500 ;
        RECT 886.8500 85.9500 888.8500 87.9500 ;
        RECT 895.0000 85.9500 897.0000 87.9500 ;
        RECT 903.1500 85.9500 905.1500 87.9500 ;
        RECT 903.1500 78.8550 905.1500 80.8550 ;
        RECT 895.0000 78.8550 897.0000 80.8550 ;
        RECT 886.8500 78.8550 888.8500 80.8550 ;
        RECT 878.7000 78.8550 880.7000 80.8550 ;
        RECT 903.1500 71.7600 905.1500 73.7600 ;
        RECT 895.0000 71.7600 897.0000 73.7600 ;
        RECT 886.8500 71.7600 888.8500 73.7600 ;
        RECT 878.7000 71.7600 880.7000 73.7600 ;
        RECT 878.7000 93.0450 880.7000 95.0450 ;
        RECT 886.8500 93.0450 888.8500 95.0450 ;
        RECT 895.0000 93.0450 897.0000 95.0450 ;
        RECT 903.1500 93.0450 905.1500 95.0450 ;
        RECT 878.7000 100.1400 880.7000 102.1400 ;
        RECT 886.8500 100.1400 888.8500 102.1400 ;
        RECT 895.0000 100.1400 897.0000 102.1400 ;
        RECT 903.1500 100.1400 905.1500 102.1400 ;
        RECT 846.1000 121.4250 848.1000 123.4250 ;
        RECT 854.2500 121.4250 856.2500 123.4250 ;
        RECT 862.4000 121.4250 864.4000 123.4250 ;
        RECT 870.5500 121.4250 872.5500 123.4250 ;
        RECT 870.5500 114.3300 872.5500 116.3300 ;
        RECT 862.4000 114.3300 864.4000 116.3300 ;
        RECT 854.2500 114.3300 856.2500 116.3300 ;
        RECT 846.1000 114.3300 848.1000 116.3300 ;
        RECT 870.5500 107.2350 872.5500 109.2350 ;
        RECT 862.4000 107.2350 864.4000 109.2350 ;
        RECT 854.2500 107.2350 856.2500 109.2350 ;
        RECT 846.1000 107.2350 848.1000 109.2350 ;
        RECT 846.1000 128.5200 848.1000 130.5200 ;
        RECT 854.2500 128.5200 856.2500 130.5200 ;
        RECT 862.4000 128.5200 864.4000 130.5200 ;
        RECT 870.5500 128.5200 872.5500 130.5200 ;
        RECT 846.1000 135.6150 848.1000 137.6150 ;
        RECT 854.2500 135.6150 856.2500 137.6150 ;
        RECT 862.4000 135.6150 864.4000 137.6150 ;
        RECT 870.5500 135.6150 872.5500 137.6150 ;
        RECT 878.7000 121.4250 880.7000 123.4250 ;
        RECT 886.8500 121.4250 888.8500 123.4250 ;
        RECT 895.0000 121.4250 897.0000 123.4250 ;
        RECT 903.1500 121.4250 905.1500 123.4250 ;
        RECT 903.1500 114.3300 905.1500 116.3300 ;
        RECT 895.0000 114.3300 897.0000 116.3300 ;
        RECT 886.8500 114.3300 888.8500 116.3300 ;
        RECT 878.7000 114.3300 880.7000 116.3300 ;
        RECT 903.1500 107.2350 905.1500 109.2350 ;
        RECT 895.0000 107.2350 897.0000 109.2350 ;
        RECT 886.8500 107.2350 888.8500 109.2350 ;
        RECT 878.7000 107.2350 880.7000 109.2350 ;
        RECT 878.7000 128.5200 880.7000 130.5200 ;
        RECT 886.8500 128.5200 888.8500 130.5200 ;
        RECT 895.0000 128.5200 897.0000 130.5200 ;
        RECT 903.1500 128.5200 905.1500 130.5200 ;
        RECT 878.7000 135.6150 880.7000 137.6150 ;
        RECT 886.8500 135.6150 888.8500 137.6150 ;
        RECT 895.0000 135.6150 897.0000 137.6150 ;
        RECT 903.1500 135.6150 905.1500 137.6150 ;
        RECT 943.9000 71.7600 945.9000 73.7600 ;
        RECT 943.9000 78.8550 945.9000 80.8550 ;
        RECT 943.9000 85.9500 945.9000 87.9500 ;
        RECT 943.9000 93.0450 945.9000 95.0450 ;
        RECT 943.9000 100.1400 945.9000 102.1400 ;
        RECT 911.3000 85.9500 913.3000 87.9500 ;
        RECT 919.4500 85.9500 921.4500 87.9500 ;
        RECT 927.6000 85.9500 929.6000 87.9500 ;
        RECT 935.7500 85.9500 937.7500 87.9500 ;
        RECT 935.7500 78.8550 937.7500 80.8550 ;
        RECT 927.6000 78.8550 929.6000 80.8550 ;
        RECT 919.4500 78.8550 921.4500 80.8550 ;
        RECT 911.3000 78.8550 913.3000 80.8550 ;
        RECT 935.7500 71.7600 937.7500 73.7600 ;
        RECT 927.6000 71.7600 929.6000 73.7600 ;
        RECT 919.4500 71.7600 921.4500 73.7600 ;
        RECT 911.3000 71.7600 913.3000 73.7600 ;
        RECT 911.3000 93.0450 913.3000 95.0450 ;
        RECT 919.4500 93.0450 921.4500 95.0450 ;
        RECT 927.6000 93.0450 929.6000 95.0450 ;
        RECT 935.7500 93.0450 937.7500 95.0450 ;
        RECT 911.3000 100.1400 913.3000 102.1400 ;
        RECT 919.4500 100.1400 921.4500 102.1400 ;
        RECT 927.6000 100.1400 929.6000 102.1400 ;
        RECT 935.7500 100.1400 937.7500 102.1400 ;
        RECT 952.0500 85.9500 954.0500 87.9500 ;
        RECT 960.2000 85.9500 962.2000 87.9500 ;
        RECT 968.3500 85.9500 970.3500 87.9500 ;
        RECT 976.5000 85.9500 978.5000 87.9500 ;
        RECT 976.5000 78.8550 978.5000 80.8550 ;
        RECT 968.3500 78.8550 970.3500 80.8550 ;
        RECT 960.2000 78.8550 962.2000 80.8550 ;
        RECT 952.0500 78.8550 954.0500 80.8550 ;
        RECT 976.5000 71.7600 978.5000 73.7600 ;
        RECT 968.3500 71.7600 970.3500 73.7600 ;
        RECT 960.2000 71.7600 962.2000 73.7600 ;
        RECT 952.0500 71.7600 954.0500 73.7600 ;
        RECT 952.0500 93.0450 954.0500 95.0450 ;
        RECT 960.2000 93.0450 962.2000 95.0450 ;
        RECT 968.3500 93.0450 970.3500 95.0450 ;
        RECT 976.5000 93.0450 978.5000 95.0450 ;
        RECT 952.0500 100.1400 954.0500 102.1400 ;
        RECT 960.2000 100.1400 962.2000 102.1400 ;
        RECT 968.3500 100.1400 970.3500 102.1400 ;
        RECT 976.5000 100.1400 978.5000 102.1400 ;
        RECT 943.9000 107.2350 945.9000 109.2350 ;
        RECT 943.9000 114.3300 945.9000 116.3300 ;
        RECT 943.9000 121.4250 945.9000 123.4250 ;
        RECT 943.9000 128.5200 945.9000 130.5200 ;
        RECT 943.9000 135.6150 945.9000 137.6150 ;
        RECT 911.3000 121.4250 913.3000 123.4250 ;
        RECT 919.4500 121.4250 921.4500 123.4250 ;
        RECT 927.6000 121.4250 929.6000 123.4250 ;
        RECT 935.7500 121.4250 937.7500 123.4250 ;
        RECT 935.7500 114.3300 937.7500 116.3300 ;
        RECT 927.6000 114.3300 929.6000 116.3300 ;
        RECT 919.4500 114.3300 921.4500 116.3300 ;
        RECT 911.3000 114.3300 913.3000 116.3300 ;
        RECT 935.7500 107.2350 937.7500 109.2350 ;
        RECT 927.6000 107.2350 929.6000 109.2350 ;
        RECT 919.4500 107.2350 921.4500 109.2350 ;
        RECT 911.3000 107.2350 913.3000 109.2350 ;
        RECT 911.3000 128.5200 913.3000 130.5200 ;
        RECT 919.4500 128.5200 921.4500 130.5200 ;
        RECT 927.6000 128.5200 929.6000 130.5200 ;
        RECT 935.7500 128.5200 937.7500 130.5200 ;
        RECT 911.3000 135.6150 913.3000 137.6150 ;
        RECT 919.4500 135.6150 921.4500 137.6150 ;
        RECT 927.6000 135.6150 929.6000 137.6150 ;
        RECT 935.7500 135.6150 937.7500 137.6150 ;
        RECT 952.0500 121.4250 954.0500 123.4250 ;
        RECT 960.2000 121.4250 962.2000 123.4250 ;
        RECT 968.3500 121.4250 970.3500 123.4250 ;
        RECT 976.5000 121.4250 978.5000 123.4250 ;
        RECT 976.5000 114.3300 978.5000 116.3300 ;
        RECT 968.3500 114.3300 970.3500 116.3300 ;
        RECT 960.2000 114.3300 962.2000 116.3300 ;
        RECT 952.0500 114.3300 954.0500 116.3300 ;
        RECT 976.5000 107.2350 978.5000 109.2350 ;
        RECT 968.3500 107.2350 970.3500 109.2350 ;
        RECT 960.2000 107.2350 962.2000 109.2350 ;
        RECT 952.0500 107.2350 954.0500 109.2350 ;
        RECT 952.0500 128.5200 954.0500 130.5200 ;
        RECT 960.2000 128.5200 962.2000 130.5200 ;
        RECT 968.3500 128.5200 970.3500 130.5200 ;
        RECT 976.5000 128.5200 978.5000 130.5200 ;
        RECT 952.0500 135.6150 954.0500 137.6150 ;
        RECT 960.2000 135.6150 962.2000 137.6150 ;
        RECT 968.3500 135.6150 970.3500 137.6150 ;
        RECT 976.5000 135.6150 978.5000 137.6150 ;
        RECT 1049.8500 64.6650 1051.8500 66.6650 ;
        RECT 984.6500 64.6650 986.6500 66.6650 ;
        RECT 992.8000 64.6650 994.8000 66.6650 ;
        RECT 1000.9500 64.6650 1002.9500 66.6650 ;
        RECT 1009.1000 64.6650 1011.1000 66.6650 ;
        RECT 1017.2500 64.6650 1019.2500 66.6650 ;
        RECT 1025.4000 64.6650 1027.4000 66.6650 ;
        RECT 1033.5500 64.6650 1035.5500 66.6650 ;
        RECT 1041.7000 64.6650 1043.7000 66.6650 ;
        RECT 1112.0000 15.0000 1114.0000 17.0000 ;
        RECT 1112.0000 22.0950 1114.0000 24.0950 ;
        RECT 1112.0000 29.1900 1114.0000 31.1900 ;
        RECT 1074.0000 44.0000 1076.0000 45.3800 ;
        RECT 1074.0000 50.4750 1076.0000 52.4750 ;
        RECT 1058.0000 64.6650 1060.0000 66.6650 ;
        RECT 1074.0000 57.5700 1076.0000 59.5700 ;
        RECT 1074.0000 64.6650 1076.0000 66.6650 ;
        RECT 1112.0000 43.3800 1114.0000 45.3800 ;
        RECT 1112.0000 36.2850 1114.0000 38.2850 ;
        RECT 1112.0000 50.4750 1114.0000 52.4750 ;
        RECT 1112.0000 57.5700 1114.0000 59.5700 ;
        RECT 1112.0000 64.6650 1114.0000 66.6650 ;
        RECT 1049.8500 71.7600 1051.8500 73.7600 ;
        RECT 1049.8500 78.8550 1051.8500 80.8550 ;
        RECT 1049.8500 85.9500 1051.8500 87.9500 ;
        RECT 1049.8500 93.0450 1051.8500 95.0450 ;
        RECT 1049.8500 100.1400 1051.8500 102.1400 ;
        RECT 1049.8500 107.2350 1051.8500 109.2350 ;
        RECT 1049.8500 114.3300 1051.8500 116.3300 ;
        RECT 1049.8500 121.4250 1051.8500 123.4250 ;
        RECT 1049.8500 128.5200 1051.8500 130.5200 ;
        RECT 1049.8500 135.6150 1051.8500 137.6150 ;
        RECT 984.6500 85.9500 986.6500 87.9500 ;
        RECT 992.8000 85.9500 994.8000 87.9500 ;
        RECT 1000.9500 85.9500 1002.9500 87.9500 ;
        RECT 1009.1000 85.9500 1011.1000 87.9500 ;
        RECT 1009.1000 78.8550 1011.1000 80.8550 ;
        RECT 1000.9500 78.8550 1002.9500 80.8550 ;
        RECT 992.8000 78.8550 994.8000 80.8550 ;
        RECT 984.6500 78.8550 986.6500 80.8550 ;
        RECT 1009.1000 71.7600 1011.1000 73.7600 ;
        RECT 1000.9500 71.7600 1002.9500 73.7600 ;
        RECT 992.8000 71.7600 994.8000 73.7600 ;
        RECT 984.6500 71.7600 986.6500 73.7600 ;
        RECT 984.6500 93.0450 986.6500 95.0450 ;
        RECT 992.8000 93.0450 994.8000 95.0450 ;
        RECT 1000.9500 93.0450 1002.9500 95.0450 ;
        RECT 1009.1000 93.0450 1011.1000 95.0450 ;
        RECT 984.6500 100.1400 986.6500 102.1400 ;
        RECT 992.8000 100.1400 994.8000 102.1400 ;
        RECT 1000.9500 100.1400 1002.9500 102.1400 ;
        RECT 1009.1000 100.1400 1011.1000 102.1400 ;
        RECT 1017.2500 85.9500 1019.2500 87.9500 ;
        RECT 1025.4000 85.9500 1027.4000 87.9500 ;
        RECT 1033.5500 85.9500 1035.5500 87.9500 ;
        RECT 1041.7000 85.9500 1043.7000 87.9500 ;
        RECT 1041.7000 78.8550 1043.7000 80.8550 ;
        RECT 1033.5500 78.8550 1035.5500 80.8550 ;
        RECT 1025.4000 78.8550 1027.4000 80.8550 ;
        RECT 1017.2500 78.8550 1019.2500 80.8550 ;
        RECT 1041.7000 71.7600 1043.7000 73.7600 ;
        RECT 1033.5500 71.7600 1035.5500 73.7600 ;
        RECT 1025.4000 71.7600 1027.4000 73.7600 ;
        RECT 1017.2500 71.7600 1019.2500 73.7600 ;
        RECT 1017.2500 93.0450 1019.2500 95.0450 ;
        RECT 1025.4000 93.0450 1027.4000 95.0450 ;
        RECT 1033.5500 93.0450 1035.5500 95.0450 ;
        RECT 1041.7000 93.0450 1043.7000 95.0450 ;
        RECT 1017.2500 100.1400 1019.2500 102.1400 ;
        RECT 1025.4000 100.1400 1027.4000 102.1400 ;
        RECT 1033.5500 100.1400 1035.5500 102.1400 ;
        RECT 1041.7000 100.1400 1043.7000 102.1400 ;
        RECT 984.6500 121.4250 986.6500 123.4250 ;
        RECT 992.8000 121.4250 994.8000 123.4250 ;
        RECT 1000.9500 121.4250 1002.9500 123.4250 ;
        RECT 1009.1000 121.4250 1011.1000 123.4250 ;
        RECT 1009.1000 114.3300 1011.1000 116.3300 ;
        RECT 1000.9500 114.3300 1002.9500 116.3300 ;
        RECT 992.8000 114.3300 994.8000 116.3300 ;
        RECT 984.6500 114.3300 986.6500 116.3300 ;
        RECT 1009.1000 107.2350 1011.1000 109.2350 ;
        RECT 1000.9500 107.2350 1002.9500 109.2350 ;
        RECT 992.8000 107.2350 994.8000 109.2350 ;
        RECT 984.6500 107.2350 986.6500 109.2350 ;
        RECT 984.6500 128.5200 986.6500 130.5200 ;
        RECT 992.8000 128.5200 994.8000 130.5200 ;
        RECT 1000.9500 128.5200 1002.9500 130.5200 ;
        RECT 1009.1000 128.5200 1011.1000 130.5200 ;
        RECT 984.6500 135.6150 986.6500 137.6150 ;
        RECT 992.8000 135.6150 994.8000 137.6150 ;
        RECT 1000.9500 135.6150 1002.9500 137.6150 ;
        RECT 1009.1000 135.6150 1011.1000 137.6150 ;
        RECT 1017.2500 121.4250 1019.2500 123.4250 ;
        RECT 1025.4000 121.4250 1027.4000 123.4250 ;
        RECT 1033.5500 121.4250 1035.5500 123.4250 ;
        RECT 1041.7000 121.4250 1043.7000 123.4250 ;
        RECT 1041.7000 114.3300 1043.7000 116.3300 ;
        RECT 1033.5500 114.3300 1035.5500 116.3300 ;
        RECT 1025.4000 114.3300 1027.4000 116.3300 ;
        RECT 1017.2500 114.3300 1019.2500 116.3300 ;
        RECT 1041.7000 107.2350 1043.7000 109.2350 ;
        RECT 1033.5500 107.2350 1035.5500 109.2350 ;
        RECT 1025.4000 107.2350 1027.4000 109.2350 ;
        RECT 1017.2500 107.2350 1019.2500 109.2350 ;
        RECT 1017.2500 128.5200 1019.2500 130.5200 ;
        RECT 1025.4000 128.5200 1027.4000 130.5200 ;
        RECT 1033.5500 128.5200 1035.5500 130.5200 ;
        RECT 1041.7000 128.5200 1043.7000 130.5200 ;
        RECT 1017.2500 135.6150 1019.2500 137.6150 ;
        RECT 1025.4000 135.6150 1027.4000 137.6150 ;
        RECT 1033.5500 135.6150 1035.5500 137.6150 ;
        RECT 1041.7000 135.6150 1043.7000 137.6150 ;
        RECT 1074.0000 85.9500 1076.0000 87.9500 ;
        RECT 1058.0000 85.9500 1060.0000 87.9500 ;
        RECT 1058.0000 78.8550 1060.0000 80.8550 ;
        RECT 1058.0000 71.7600 1060.0000 73.7600 ;
        RECT 1074.0000 78.8550 1076.0000 80.8550 ;
        RECT 1074.0000 71.7600 1076.0000 73.7600 ;
        RECT 1058.0000 100.1400 1060.0000 102.1400 ;
        RECT 1058.0000 93.0450 1060.0000 95.0450 ;
        RECT 1074.0000 93.0450 1076.0000 95.0450 ;
        RECT 1074.0000 100.1400 1076.0000 102.1400 ;
        RECT 1112.0000 85.9500 1114.0000 87.9500 ;
        RECT 1112.0000 71.7600 1114.0000 73.7600 ;
        RECT 1112.0000 78.8550 1114.0000 80.8550 ;
        RECT 1112.0000 93.0450 1114.0000 95.0450 ;
        RECT 1112.0000 100.1400 1114.0000 102.1400 ;
        RECT 1074.0000 121.4250 1076.0000 123.4250 ;
        RECT 1058.0000 121.4250 1060.0000 123.4250 ;
        RECT 1058.0000 114.3300 1060.0000 116.3300 ;
        RECT 1058.0000 107.2350 1060.0000 109.2350 ;
        RECT 1074.0000 107.2350 1076.0000 109.2350 ;
        RECT 1074.0000 114.3300 1076.0000 116.3300 ;
        RECT 1058.0000 135.6150 1060.0000 137.6150 ;
        RECT 1058.0000 128.5200 1060.0000 130.5200 ;
        RECT 1074.0000 128.5200 1076.0000 130.5200 ;
        RECT 1074.0000 135.6150 1076.0000 137.6150 ;
        RECT 1112.0000 121.4250 1114.0000 123.4250 ;
        RECT 1112.0000 107.2350 1114.0000 109.2350 ;
        RECT 1112.0000 114.3300 1114.0000 116.3300 ;
        RECT 1112.0000 128.5200 1114.0000 130.5200 ;
        RECT 1112.0000 135.6150 1114.0000 137.6150 ;
        RECT 846.1000 156.9000 848.1000 158.9000 ;
        RECT 854.2500 156.9000 856.2500 158.9000 ;
        RECT 862.4000 156.9000 864.4000 158.9000 ;
        RECT 870.5500 156.9000 872.5500 158.9000 ;
        RECT 870.5500 149.8050 872.5500 151.8050 ;
        RECT 862.4000 149.8050 864.4000 151.8050 ;
        RECT 854.2500 149.8050 856.2500 151.8050 ;
        RECT 846.1000 149.8050 848.1000 151.8050 ;
        RECT 870.5500 142.7100 872.5500 144.7100 ;
        RECT 862.4000 142.7100 864.4000 144.7100 ;
        RECT 854.2500 142.7100 856.2500 144.7100 ;
        RECT 846.1000 142.7100 848.1000 144.7100 ;
        RECT 846.1000 163.9950 848.1000 165.9950 ;
        RECT 854.2500 163.9950 856.2500 165.9950 ;
        RECT 862.4000 163.9950 864.4000 165.9950 ;
        RECT 870.5500 163.9950 872.5500 165.9950 ;
        RECT 846.1000 171.0900 848.1000 173.0900 ;
        RECT 854.2500 171.0900 856.2500 173.0900 ;
        RECT 862.4000 171.0900 864.4000 173.0900 ;
        RECT 870.5500 171.0900 872.5500 173.0900 ;
        RECT 878.7000 156.9000 880.7000 158.9000 ;
        RECT 886.8500 156.9000 888.8500 158.9000 ;
        RECT 895.0000 156.9000 897.0000 158.9000 ;
        RECT 903.1500 156.9000 905.1500 158.9000 ;
        RECT 903.1500 149.8050 905.1500 151.8050 ;
        RECT 895.0000 149.8050 897.0000 151.8050 ;
        RECT 886.8500 149.8050 888.8500 151.8050 ;
        RECT 878.7000 149.8050 880.7000 151.8050 ;
        RECT 903.1500 142.7100 905.1500 144.7100 ;
        RECT 895.0000 142.7100 897.0000 144.7100 ;
        RECT 886.8500 142.7100 888.8500 144.7100 ;
        RECT 878.7000 142.7100 880.7000 144.7100 ;
        RECT 878.7000 163.9950 880.7000 165.9950 ;
        RECT 886.8500 163.9950 888.8500 165.9950 ;
        RECT 895.0000 163.9950 897.0000 165.9950 ;
        RECT 903.1500 163.9950 905.1500 165.9950 ;
        RECT 878.7000 171.0900 880.7000 173.0900 ;
        RECT 886.8500 171.0900 888.8500 173.0900 ;
        RECT 895.0000 171.0900 897.0000 173.0900 ;
        RECT 903.1500 171.0900 905.1500 173.0900 ;
        RECT 846.1000 192.3750 848.1000 194.3750 ;
        RECT 854.2500 192.3750 856.2500 194.3750 ;
        RECT 862.4000 192.3750 864.4000 194.3750 ;
        RECT 870.5500 192.3750 872.5500 194.3750 ;
        RECT 870.5500 185.2800 872.5500 187.2800 ;
        RECT 862.4000 185.2800 864.4000 187.2800 ;
        RECT 854.2500 185.2800 856.2500 187.2800 ;
        RECT 846.1000 185.2800 848.1000 187.2800 ;
        RECT 870.5500 178.1850 872.5500 180.1850 ;
        RECT 862.4000 178.1850 864.4000 180.1850 ;
        RECT 854.2500 178.1850 856.2500 180.1850 ;
        RECT 846.1000 178.1850 848.1000 180.1850 ;
        RECT 846.1000 199.4700 848.1000 201.4700 ;
        RECT 854.2500 199.4700 856.2500 201.4700 ;
        RECT 862.4000 199.4700 864.4000 201.4700 ;
        RECT 870.5500 199.4700 872.5500 201.4700 ;
        RECT 846.1000 206.5650 848.1000 208.5650 ;
        RECT 854.2500 206.5650 856.2500 208.5650 ;
        RECT 862.4000 206.5650 864.4000 208.5650 ;
        RECT 870.5500 206.5650 872.5500 208.5650 ;
        RECT 878.7000 192.3750 880.7000 194.3750 ;
        RECT 886.8500 192.3750 888.8500 194.3750 ;
        RECT 895.0000 192.3750 897.0000 194.3750 ;
        RECT 903.1500 192.3750 905.1500 194.3750 ;
        RECT 903.1500 185.2800 905.1500 187.2800 ;
        RECT 895.0000 185.2800 897.0000 187.2800 ;
        RECT 886.8500 185.2800 888.8500 187.2800 ;
        RECT 878.7000 185.2800 880.7000 187.2800 ;
        RECT 903.1500 178.1850 905.1500 180.1850 ;
        RECT 895.0000 178.1850 897.0000 180.1850 ;
        RECT 886.8500 178.1850 888.8500 180.1850 ;
        RECT 878.7000 178.1850 880.7000 180.1850 ;
        RECT 878.7000 199.4700 880.7000 201.4700 ;
        RECT 886.8500 199.4700 888.8500 201.4700 ;
        RECT 895.0000 199.4700 897.0000 201.4700 ;
        RECT 903.1500 199.4700 905.1500 201.4700 ;
        RECT 878.7000 206.5650 880.7000 208.5650 ;
        RECT 886.8500 206.5650 888.8500 208.5650 ;
        RECT 895.0000 206.5650 897.0000 208.5650 ;
        RECT 903.1500 206.5650 905.1500 208.5650 ;
        RECT 943.9000 142.7100 945.9000 144.7100 ;
        RECT 943.9000 149.8050 945.9000 151.8050 ;
        RECT 943.9000 156.9000 945.9000 158.9000 ;
        RECT 943.9000 163.9950 945.9000 165.9950 ;
        RECT 943.9000 171.0900 945.9000 173.0900 ;
        RECT 911.3000 156.9000 913.3000 158.9000 ;
        RECT 919.4500 156.9000 921.4500 158.9000 ;
        RECT 927.6000 156.9000 929.6000 158.9000 ;
        RECT 935.7500 156.9000 937.7500 158.9000 ;
        RECT 935.7500 149.8050 937.7500 151.8050 ;
        RECT 927.6000 149.8050 929.6000 151.8050 ;
        RECT 919.4500 149.8050 921.4500 151.8050 ;
        RECT 911.3000 149.8050 913.3000 151.8050 ;
        RECT 935.7500 142.7100 937.7500 144.7100 ;
        RECT 927.6000 142.7100 929.6000 144.7100 ;
        RECT 919.4500 142.7100 921.4500 144.7100 ;
        RECT 911.3000 142.7100 913.3000 144.7100 ;
        RECT 911.3000 163.9950 913.3000 165.9950 ;
        RECT 919.4500 163.9950 921.4500 165.9950 ;
        RECT 927.6000 163.9950 929.6000 165.9950 ;
        RECT 935.7500 163.9950 937.7500 165.9950 ;
        RECT 911.3000 171.0900 913.3000 173.0900 ;
        RECT 919.4500 171.0900 921.4500 173.0900 ;
        RECT 927.6000 171.0900 929.6000 173.0900 ;
        RECT 935.7500 171.0900 937.7500 173.0900 ;
        RECT 952.0500 156.9000 954.0500 158.9000 ;
        RECT 960.2000 156.9000 962.2000 158.9000 ;
        RECT 968.3500 156.9000 970.3500 158.9000 ;
        RECT 976.5000 156.9000 978.5000 158.9000 ;
        RECT 976.5000 149.8050 978.5000 151.8050 ;
        RECT 968.3500 149.8050 970.3500 151.8050 ;
        RECT 960.2000 149.8050 962.2000 151.8050 ;
        RECT 952.0500 149.8050 954.0500 151.8050 ;
        RECT 976.5000 142.7100 978.5000 144.7100 ;
        RECT 968.3500 142.7100 970.3500 144.7100 ;
        RECT 960.2000 142.7100 962.2000 144.7100 ;
        RECT 952.0500 142.7100 954.0500 144.7100 ;
        RECT 952.0500 163.9950 954.0500 165.9950 ;
        RECT 960.2000 163.9950 962.2000 165.9950 ;
        RECT 968.3500 163.9950 970.3500 165.9950 ;
        RECT 976.5000 163.9950 978.5000 165.9950 ;
        RECT 952.0500 171.0900 954.0500 173.0900 ;
        RECT 960.2000 171.0900 962.2000 173.0900 ;
        RECT 968.3500 171.0900 970.3500 173.0900 ;
        RECT 976.5000 171.0900 978.5000 173.0900 ;
        RECT 943.9000 178.1850 945.9000 180.1850 ;
        RECT 943.9000 185.2800 945.9000 187.2800 ;
        RECT 943.9000 192.3750 945.9000 194.3750 ;
        RECT 943.9000 199.4700 945.9000 201.4700 ;
        RECT 943.9000 206.5650 945.9000 208.5650 ;
        RECT 911.3000 192.3750 913.3000 194.3750 ;
        RECT 919.4500 192.3750 921.4500 194.3750 ;
        RECT 927.6000 192.3750 929.6000 194.3750 ;
        RECT 935.7500 192.3750 937.7500 194.3750 ;
        RECT 935.7500 185.2800 937.7500 187.2800 ;
        RECT 927.6000 185.2800 929.6000 187.2800 ;
        RECT 919.4500 185.2800 921.4500 187.2800 ;
        RECT 911.3000 185.2800 913.3000 187.2800 ;
        RECT 935.7500 178.1850 937.7500 180.1850 ;
        RECT 927.6000 178.1850 929.6000 180.1850 ;
        RECT 919.4500 178.1850 921.4500 180.1850 ;
        RECT 911.3000 178.1850 913.3000 180.1850 ;
        RECT 911.3000 199.4700 913.3000 201.4700 ;
        RECT 919.4500 199.4700 921.4500 201.4700 ;
        RECT 927.6000 199.4700 929.6000 201.4700 ;
        RECT 935.7500 199.4700 937.7500 201.4700 ;
        RECT 911.3000 206.5650 913.3000 208.5650 ;
        RECT 919.4500 206.5650 921.4500 208.5650 ;
        RECT 927.6000 206.5650 929.6000 208.5650 ;
        RECT 935.7500 206.5650 937.7500 208.5650 ;
        RECT 952.0500 192.3750 954.0500 194.3750 ;
        RECT 960.2000 192.3750 962.2000 194.3750 ;
        RECT 968.3500 192.3750 970.3500 194.3750 ;
        RECT 976.5000 192.3750 978.5000 194.3750 ;
        RECT 976.5000 185.2800 978.5000 187.2800 ;
        RECT 968.3500 185.2800 970.3500 187.2800 ;
        RECT 960.2000 185.2800 962.2000 187.2800 ;
        RECT 952.0500 185.2800 954.0500 187.2800 ;
        RECT 976.5000 178.1850 978.5000 180.1850 ;
        RECT 968.3500 178.1850 970.3500 180.1850 ;
        RECT 960.2000 178.1850 962.2000 180.1850 ;
        RECT 952.0500 178.1850 954.0500 180.1850 ;
        RECT 952.0500 199.4700 954.0500 201.4700 ;
        RECT 960.2000 199.4700 962.2000 201.4700 ;
        RECT 968.3500 199.4700 970.3500 201.4700 ;
        RECT 976.5000 199.4700 978.5000 201.4700 ;
        RECT 952.0500 206.5650 954.0500 208.5650 ;
        RECT 960.2000 206.5650 962.2000 208.5650 ;
        RECT 968.3500 206.5650 970.3500 208.5650 ;
        RECT 976.5000 206.5650 978.5000 208.5650 ;
        RECT 870.5500 220.7550 872.5500 222.7550 ;
        RECT 862.4000 220.7550 864.4000 222.7550 ;
        RECT 854.2500 220.7550 856.2500 222.7550 ;
        RECT 846.1000 220.7550 848.1000 222.7550 ;
        RECT 870.5500 213.6600 872.5500 215.6600 ;
        RECT 862.4000 213.6600 864.4000 215.6600 ;
        RECT 854.2500 213.6600 856.2500 215.6600 ;
        RECT 846.1000 213.6600 848.1000 215.6600 ;
        RECT 854.2500 227.8500 856.2500 229.8500 ;
        RECT 846.1000 227.8500 848.1000 229.8500 ;
        RECT 862.4000 227.8500 864.4000 229.8500 ;
        RECT 870.5500 227.8500 872.5500 229.8500 ;
        RECT 846.1000 234.9450 848.1000 236.9450 ;
        RECT 854.2500 234.9450 856.2500 236.9450 ;
        RECT 862.4000 234.9450 864.4000 236.9450 ;
        RECT 870.5500 234.9450 872.5500 236.9450 ;
        RECT 846.1000 242.0400 848.1000 244.0400 ;
        RECT 854.2500 242.0400 856.2500 244.0400 ;
        RECT 862.4000 242.0400 864.4000 244.0400 ;
        RECT 870.5500 242.0400 872.5500 244.0400 ;
        RECT 903.1500 220.7550 905.1500 222.7550 ;
        RECT 895.0000 220.7550 897.0000 222.7550 ;
        RECT 886.8500 220.7550 888.8500 222.7550 ;
        RECT 878.7000 220.7550 880.7000 222.7550 ;
        RECT 903.1500 213.6600 905.1500 215.6600 ;
        RECT 895.0000 213.6600 897.0000 215.6600 ;
        RECT 886.8500 213.6600 888.8500 215.6600 ;
        RECT 878.7000 213.6600 880.7000 215.6600 ;
        RECT 886.8500 227.8500 888.8500 229.8500 ;
        RECT 878.7000 227.8500 880.7000 229.8500 ;
        RECT 895.0000 227.8500 897.0000 229.8500 ;
        RECT 903.1500 227.8500 905.1500 229.8500 ;
        RECT 878.7000 234.9450 880.7000 236.9450 ;
        RECT 886.8500 234.9450 888.8500 236.9450 ;
        RECT 895.0000 234.9450 897.0000 236.9450 ;
        RECT 903.1500 234.9450 905.1500 236.9450 ;
        RECT 878.7000 242.0400 880.7000 244.0400 ;
        RECT 886.8500 242.0400 888.8500 244.0400 ;
        RECT 895.0000 242.0400 897.0000 244.0400 ;
        RECT 903.1500 242.0400 905.1500 244.0400 ;
        RECT 870.5500 256.2300 872.5500 258.2300 ;
        RECT 862.4000 256.2300 864.4000 258.2300 ;
        RECT 854.2500 256.2300 856.2500 258.2300 ;
        RECT 846.1000 256.2300 848.1000 258.2300 ;
        RECT 870.5500 249.1350 872.5500 251.1350 ;
        RECT 862.4000 249.1350 864.4000 251.1350 ;
        RECT 854.2500 249.1350 856.2500 251.1350 ;
        RECT 846.1000 249.1350 848.1000 251.1350 ;
        RECT 854.2500 263.3250 856.2500 265.3250 ;
        RECT 846.1000 263.3250 848.1000 265.3250 ;
        RECT 862.4000 263.3250 864.4000 265.3250 ;
        RECT 870.5500 263.3250 872.5500 265.3250 ;
        RECT 846.1000 270.4200 848.1000 272.4200 ;
        RECT 854.2500 270.4200 856.2500 272.4200 ;
        RECT 862.4000 270.4200 864.4000 272.4200 ;
        RECT 870.5500 270.4200 872.5500 272.4200 ;
        RECT 846.1000 277.5150 848.1000 279.5150 ;
        RECT 854.2500 277.5150 856.2500 279.5150 ;
        RECT 862.4000 277.5150 864.4000 279.5150 ;
        RECT 870.5500 277.5150 872.5500 279.5150 ;
        RECT 903.1500 256.2300 905.1500 258.2300 ;
        RECT 895.0000 256.2300 897.0000 258.2300 ;
        RECT 886.8500 256.2300 888.8500 258.2300 ;
        RECT 878.7000 256.2300 880.7000 258.2300 ;
        RECT 903.1500 249.1350 905.1500 251.1350 ;
        RECT 895.0000 249.1350 897.0000 251.1350 ;
        RECT 886.8500 249.1350 888.8500 251.1350 ;
        RECT 878.7000 249.1350 880.7000 251.1350 ;
        RECT 886.8500 263.3250 888.8500 265.3250 ;
        RECT 878.7000 263.3250 880.7000 265.3250 ;
        RECT 895.0000 263.3250 897.0000 265.3250 ;
        RECT 903.1500 263.3250 905.1500 265.3250 ;
        RECT 878.7000 270.4200 880.7000 272.4200 ;
        RECT 886.8500 270.4200 888.8500 272.4200 ;
        RECT 895.0000 270.4200 897.0000 272.4200 ;
        RECT 903.1500 270.4200 905.1500 272.4200 ;
        RECT 878.7000 277.5150 880.7000 279.5150 ;
        RECT 886.8500 277.5150 888.8500 279.5150 ;
        RECT 895.0000 277.5150 897.0000 279.5150 ;
        RECT 903.1500 277.5150 905.1500 279.5150 ;
        RECT 943.9000 213.6600 945.9000 215.6600 ;
        RECT 943.9000 220.7550 945.9000 222.7550 ;
        RECT 943.9000 227.8500 945.9000 229.8500 ;
        RECT 943.9000 234.9450 945.9000 236.9450 ;
        RECT 943.9000 242.0400 945.9000 244.0400 ;
        RECT 935.7500 220.7550 937.7500 222.7550 ;
        RECT 927.6000 220.7550 929.6000 222.7550 ;
        RECT 919.4500 220.7550 921.4500 222.7550 ;
        RECT 911.3000 220.7550 913.3000 222.7550 ;
        RECT 935.7500 213.6600 937.7500 215.6600 ;
        RECT 927.6000 213.6600 929.6000 215.6600 ;
        RECT 919.4500 213.6600 921.4500 215.6600 ;
        RECT 911.3000 213.6600 913.3000 215.6600 ;
        RECT 919.4500 227.8500 921.4500 229.8500 ;
        RECT 911.3000 227.8500 913.3000 229.8500 ;
        RECT 927.6000 227.8500 929.6000 229.8500 ;
        RECT 935.7500 227.8500 937.7500 229.8500 ;
        RECT 911.3000 234.9450 913.3000 236.9450 ;
        RECT 919.4500 234.9450 921.4500 236.9450 ;
        RECT 927.6000 234.9450 929.6000 236.9450 ;
        RECT 935.7500 234.9450 937.7500 236.9450 ;
        RECT 911.3000 242.0400 913.3000 244.0400 ;
        RECT 919.4500 242.0400 921.4500 244.0400 ;
        RECT 927.6000 242.0400 929.6000 244.0400 ;
        RECT 935.7500 242.0400 937.7500 244.0400 ;
        RECT 976.5000 220.7550 978.5000 222.7550 ;
        RECT 968.3500 220.7550 970.3500 222.7550 ;
        RECT 960.2000 220.7550 962.2000 222.7550 ;
        RECT 952.0500 220.7550 954.0500 222.7550 ;
        RECT 976.5000 213.6600 978.5000 215.6600 ;
        RECT 968.3500 213.6600 970.3500 215.6600 ;
        RECT 960.2000 213.6600 962.2000 215.6600 ;
        RECT 952.0500 213.6600 954.0500 215.6600 ;
        RECT 960.2000 227.8500 962.2000 229.8500 ;
        RECT 952.0500 227.8500 954.0500 229.8500 ;
        RECT 968.3500 227.8500 970.3500 229.8500 ;
        RECT 976.5000 227.8500 978.5000 229.8500 ;
        RECT 952.0500 234.9450 954.0500 236.9450 ;
        RECT 960.2000 234.9450 962.2000 236.9450 ;
        RECT 968.3500 234.9450 970.3500 236.9450 ;
        RECT 976.5000 234.9450 978.5000 236.9450 ;
        RECT 952.0500 242.0400 954.0500 244.0400 ;
        RECT 960.2000 242.0400 962.2000 244.0400 ;
        RECT 968.3500 242.0400 970.3500 244.0400 ;
        RECT 976.5000 242.0400 978.5000 244.0400 ;
        RECT 943.9000 249.1350 945.9000 251.1350 ;
        RECT 943.9000 256.2300 945.9000 258.2300 ;
        RECT 943.9000 263.3250 945.9000 265.3250 ;
        RECT 943.9000 270.4200 945.9000 272.4200 ;
        RECT 943.9000 277.5150 945.9000 279.5150 ;
        RECT 935.7500 256.2300 937.7500 258.2300 ;
        RECT 927.6000 256.2300 929.6000 258.2300 ;
        RECT 919.4500 256.2300 921.4500 258.2300 ;
        RECT 911.3000 256.2300 913.3000 258.2300 ;
        RECT 935.7500 249.1350 937.7500 251.1350 ;
        RECT 927.6000 249.1350 929.6000 251.1350 ;
        RECT 919.4500 249.1350 921.4500 251.1350 ;
        RECT 911.3000 249.1350 913.3000 251.1350 ;
        RECT 919.4500 263.3250 921.4500 265.3250 ;
        RECT 911.3000 263.3250 913.3000 265.3250 ;
        RECT 927.6000 263.3250 929.6000 265.3250 ;
        RECT 935.7500 263.3250 937.7500 265.3250 ;
        RECT 911.3000 270.4200 913.3000 272.4200 ;
        RECT 919.4500 270.4200 921.4500 272.4200 ;
        RECT 927.6000 270.4200 929.6000 272.4200 ;
        RECT 935.7500 270.4200 937.7500 272.4200 ;
        RECT 911.3000 277.5150 913.3000 279.5150 ;
        RECT 919.4500 277.5150 921.4500 279.5150 ;
        RECT 927.6000 277.5150 929.6000 279.5150 ;
        RECT 935.7500 277.5150 937.7500 279.5150 ;
        RECT 976.5000 256.2300 978.5000 258.2300 ;
        RECT 968.3500 256.2300 970.3500 258.2300 ;
        RECT 960.2000 256.2300 962.2000 258.2300 ;
        RECT 952.0500 256.2300 954.0500 258.2300 ;
        RECT 976.5000 249.1350 978.5000 251.1350 ;
        RECT 968.3500 249.1350 970.3500 251.1350 ;
        RECT 960.2000 249.1350 962.2000 251.1350 ;
        RECT 952.0500 249.1350 954.0500 251.1350 ;
        RECT 960.2000 263.3250 962.2000 265.3250 ;
        RECT 952.0500 263.3250 954.0500 265.3250 ;
        RECT 968.3500 263.3250 970.3500 265.3250 ;
        RECT 976.5000 263.3250 978.5000 265.3250 ;
        RECT 952.0500 270.4200 954.0500 272.4200 ;
        RECT 960.2000 270.4200 962.2000 272.4200 ;
        RECT 968.3500 270.4200 970.3500 272.4200 ;
        RECT 976.5000 270.4200 978.5000 272.4200 ;
        RECT 952.0500 277.5150 954.0500 279.5150 ;
        RECT 960.2000 277.5150 962.2000 279.5150 ;
        RECT 968.3500 277.5150 970.3500 279.5150 ;
        RECT 976.5000 277.5150 978.5000 279.5150 ;
        RECT 1049.8500 142.7100 1051.8500 144.7100 ;
        RECT 1049.8500 149.8050 1051.8500 151.8050 ;
        RECT 1049.8500 156.9000 1051.8500 158.9000 ;
        RECT 1049.8500 163.9950 1051.8500 165.9950 ;
        RECT 1049.8500 171.0900 1051.8500 173.0900 ;
        RECT 1049.8500 178.1850 1051.8500 180.1850 ;
        RECT 1049.8500 185.2800 1051.8500 187.2800 ;
        RECT 1049.8500 192.3750 1051.8500 194.3750 ;
        RECT 1049.8500 199.4700 1051.8500 201.4700 ;
        RECT 1049.8500 206.5650 1051.8500 208.5650 ;
        RECT 984.6500 156.9000 986.6500 158.9000 ;
        RECT 992.8000 156.9000 994.8000 158.9000 ;
        RECT 1000.9500 156.9000 1002.9500 158.9000 ;
        RECT 1009.1000 156.9000 1011.1000 158.9000 ;
        RECT 1009.1000 149.8050 1011.1000 151.8050 ;
        RECT 1000.9500 149.8050 1002.9500 151.8050 ;
        RECT 992.8000 149.8050 994.8000 151.8050 ;
        RECT 984.6500 149.8050 986.6500 151.8050 ;
        RECT 1009.1000 142.7100 1011.1000 144.7100 ;
        RECT 1000.9500 142.7100 1002.9500 144.7100 ;
        RECT 992.8000 142.7100 994.8000 144.7100 ;
        RECT 984.6500 142.7100 986.6500 144.7100 ;
        RECT 984.6500 163.9950 986.6500 165.9950 ;
        RECT 992.8000 163.9950 994.8000 165.9950 ;
        RECT 1000.9500 163.9950 1002.9500 165.9950 ;
        RECT 1009.1000 163.9950 1011.1000 165.9950 ;
        RECT 984.6500 171.0900 986.6500 173.0900 ;
        RECT 992.8000 171.0900 994.8000 173.0900 ;
        RECT 1000.9500 171.0900 1002.9500 173.0900 ;
        RECT 1009.1000 171.0900 1011.1000 173.0900 ;
        RECT 1017.2500 156.9000 1019.2500 158.9000 ;
        RECT 1025.4000 156.9000 1027.4000 158.9000 ;
        RECT 1033.5500 156.9000 1035.5500 158.9000 ;
        RECT 1041.7000 156.9000 1043.7000 158.9000 ;
        RECT 1041.7000 149.8050 1043.7000 151.8050 ;
        RECT 1033.5500 149.8050 1035.5500 151.8050 ;
        RECT 1025.4000 149.8050 1027.4000 151.8050 ;
        RECT 1017.2500 149.8050 1019.2500 151.8050 ;
        RECT 1041.7000 142.7100 1043.7000 144.7100 ;
        RECT 1033.5500 142.7100 1035.5500 144.7100 ;
        RECT 1025.4000 142.7100 1027.4000 144.7100 ;
        RECT 1017.2500 142.7100 1019.2500 144.7100 ;
        RECT 1017.2500 163.9950 1019.2500 165.9950 ;
        RECT 1025.4000 163.9950 1027.4000 165.9950 ;
        RECT 1033.5500 163.9950 1035.5500 165.9950 ;
        RECT 1041.7000 163.9950 1043.7000 165.9950 ;
        RECT 1017.2500 171.0900 1019.2500 173.0900 ;
        RECT 1025.4000 171.0900 1027.4000 173.0900 ;
        RECT 1033.5500 171.0900 1035.5500 173.0900 ;
        RECT 1041.7000 171.0900 1043.7000 173.0900 ;
        RECT 984.6500 192.3750 986.6500 194.3750 ;
        RECT 992.8000 192.3750 994.8000 194.3750 ;
        RECT 1000.9500 192.3750 1002.9500 194.3750 ;
        RECT 1009.1000 192.3750 1011.1000 194.3750 ;
        RECT 1009.1000 185.2800 1011.1000 187.2800 ;
        RECT 1000.9500 185.2800 1002.9500 187.2800 ;
        RECT 992.8000 185.2800 994.8000 187.2800 ;
        RECT 984.6500 185.2800 986.6500 187.2800 ;
        RECT 1009.1000 178.1850 1011.1000 180.1850 ;
        RECT 1000.9500 178.1850 1002.9500 180.1850 ;
        RECT 992.8000 178.1850 994.8000 180.1850 ;
        RECT 984.6500 178.1850 986.6500 180.1850 ;
        RECT 984.6500 199.4700 986.6500 201.4700 ;
        RECT 992.8000 199.4700 994.8000 201.4700 ;
        RECT 1000.9500 199.4700 1002.9500 201.4700 ;
        RECT 1009.1000 199.4700 1011.1000 201.4700 ;
        RECT 984.6500 206.5650 986.6500 208.5650 ;
        RECT 992.8000 206.5650 994.8000 208.5650 ;
        RECT 1000.9500 206.5650 1002.9500 208.5650 ;
        RECT 1009.1000 206.5650 1011.1000 208.5650 ;
        RECT 1017.2500 192.3750 1019.2500 194.3750 ;
        RECT 1025.4000 192.3750 1027.4000 194.3750 ;
        RECT 1033.5500 192.3750 1035.5500 194.3750 ;
        RECT 1041.7000 192.3750 1043.7000 194.3750 ;
        RECT 1041.7000 185.2800 1043.7000 187.2800 ;
        RECT 1033.5500 185.2800 1035.5500 187.2800 ;
        RECT 1025.4000 185.2800 1027.4000 187.2800 ;
        RECT 1017.2500 185.2800 1019.2500 187.2800 ;
        RECT 1041.7000 178.1850 1043.7000 180.1850 ;
        RECT 1033.5500 178.1850 1035.5500 180.1850 ;
        RECT 1025.4000 178.1850 1027.4000 180.1850 ;
        RECT 1017.2500 178.1850 1019.2500 180.1850 ;
        RECT 1017.2500 199.4700 1019.2500 201.4700 ;
        RECT 1025.4000 199.4700 1027.4000 201.4700 ;
        RECT 1033.5500 199.4700 1035.5500 201.4700 ;
        RECT 1041.7000 199.4700 1043.7000 201.4700 ;
        RECT 1017.2500 206.5650 1019.2500 208.5650 ;
        RECT 1025.4000 206.5650 1027.4000 208.5650 ;
        RECT 1033.5500 206.5650 1035.5500 208.5650 ;
        RECT 1041.7000 206.5650 1043.7000 208.5650 ;
        RECT 1074.0000 156.9000 1076.0000 158.9000 ;
        RECT 1058.0000 156.9000 1060.0000 158.9000 ;
        RECT 1058.0000 149.8050 1060.0000 151.8050 ;
        RECT 1058.0000 142.7100 1060.0000 144.7100 ;
        RECT 1074.0000 149.8050 1076.0000 151.8050 ;
        RECT 1074.0000 142.7100 1076.0000 144.7100 ;
        RECT 1058.0000 171.0900 1060.0000 173.0900 ;
        RECT 1058.0000 163.9950 1060.0000 165.9950 ;
        RECT 1074.0000 171.0900 1076.0000 173.0900 ;
        RECT 1074.0000 163.9950 1076.0000 165.9950 ;
        RECT 1112.0000 156.9000 1114.0000 158.9000 ;
        RECT 1112.0000 142.7100 1114.0000 144.7100 ;
        RECT 1112.0000 149.8050 1114.0000 151.8050 ;
        RECT 1112.0000 163.9950 1114.0000 165.9950 ;
        RECT 1112.0000 171.0900 1114.0000 173.0900 ;
        RECT 1074.0000 192.3750 1076.0000 194.3750 ;
        RECT 1058.0000 192.3750 1060.0000 194.3750 ;
        RECT 1058.0000 185.2800 1060.0000 187.2800 ;
        RECT 1058.0000 178.1850 1060.0000 180.1850 ;
        RECT 1074.0000 178.1850 1076.0000 180.1850 ;
        RECT 1074.0000 185.2800 1076.0000 187.2800 ;
        RECT 1058.0000 206.5650 1060.0000 208.5650 ;
        RECT 1058.0000 199.4700 1060.0000 201.4700 ;
        RECT 1074.0000 199.4700 1076.0000 201.4700 ;
        RECT 1074.0000 206.5650 1076.0000 208.5650 ;
        RECT 1112.0000 192.3750 1114.0000 194.3750 ;
        RECT 1112.0000 178.1850 1114.0000 180.1850 ;
        RECT 1112.0000 185.2800 1114.0000 187.2800 ;
        RECT 1112.0000 199.4700 1114.0000 201.4700 ;
        RECT 1112.0000 206.5650 1114.0000 208.5650 ;
        RECT 1049.8500 213.6600 1051.8500 215.6600 ;
        RECT 1049.8500 220.7550 1051.8500 222.7550 ;
        RECT 1049.8500 227.8500 1051.8500 229.8500 ;
        RECT 1049.8500 234.9450 1051.8500 236.9450 ;
        RECT 1049.8500 242.0400 1051.8500 244.0400 ;
        RECT 1049.8500 249.1350 1051.8500 251.1350 ;
        RECT 1049.8500 256.2300 1051.8500 258.2300 ;
        RECT 1049.8500 263.3250 1051.8500 265.3250 ;
        RECT 1049.8500 270.4200 1051.8500 272.4200 ;
        RECT 1049.8500 277.5150 1051.8500 279.5150 ;
        RECT 1009.1000 220.7550 1011.1000 222.7550 ;
        RECT 1000.9500 220.7550 1002.9500 222.7550 ;
        RECT 992.8000 220.7550 994.8000 222.7550 ;
        RECT 984.6500 220.7550 986.6500 222.7550 ;
        RECT 1009.1000 213.6600 1011.1000 215.6600 ;
        RECT 1000.9500 213.6600 1002.9500 215.6600 ;
        RECT 992.8000 213.6600 994.8000 215.6600 ;
        RECT 984.6500 213.6600 986.6500 215.6600 ;
        RECT 992.8000 227.8500 994.8000 229.8500 ;
        RECT 984.6500 227.8500 986.6500 229.8500 ;
        RECT 1000.9500 227.8500 1002.9500 229.8500 ;
        RECT 1009.1000 227.8500 1011.1000 229.8500 ;
        RECT 984.6500 234.9450 986.6500 236.9450 ;
        RECT 992.8000 234.9450 994.8000 236.9450 ;
        RECT 1000.9500 234.9450 1002.9500 236.9450 ;
        RECT 1009.1000 234.9450 1011.1000 236.9450 ;
        RECT 984.6500 242.0400 986.6500 244.0400 ;
        RECT 992.8000 242.0400 994.8000 244.0400 ;
        RECT 1000.9500 242.0400 1002.9500 244.0400 ;
        RECT 1009.1000 242.0400 1011.1000 244.0400 ;
        RECT 1041.7000 220.7550 1043.7000 222.7550 ;
        RECT 1033.5500 220.7550 1035.5500 222.7550 ;
        RECT 1025.4000 220.7550 1027.4000 222.7550 ;
        RECT 1017.2500 220.7550 1019.2500 222.7550 ;
        RECT 1041.7000 213.6600 1043.7000 215.6600 ;
        RECT 1033.5500 213.6600 1035.5500 215.6600 ;
        RECT 1025.4000 213.6600 1027.4000 215.6600 ;
        RECT 1017.2500 213.6600 1019.2500 215.6600 ;
        RECT 1025.4000 227.8500 1027.4000 229.8500 ;
        RECT 1017.2500 227.8500 1019.2500 229.8500 ;
        RECT 1033.5500 227.8500 1035.5500 229.8500 ;
        RECT 1041.7000 227.8500 1043.7000 229.8500 ;
        RECT 1017.2500 234.9450 1019.2500 236.9450 ;
        RECT 1025.4000 234.9450 1027.4000 236.9450 ;
        RECT 1033.5500 234.9450 1035.5500 236.9450 ;
        RECT 1041.7000 234.9450 1043.7000 236.9450 ;
        RECT 1017.2500 242.0400 1019.2500 244.0400 ;
        RECT 1025.4000 242.0400 1027.4000 244.0400 ;
        RECT 1033.5500 242.0400 1035.5500 244.0400 ;
        RECT 1041.7000 242.0400 1043.7000 244.0400 ;
        RECT 1009.1000 256.2300 1011.1000 258.2300 ;
        RECT 1000.9500 256.2300 1002.9500 258.2300 ;
        RECT 992.8000 256.2300 994.8000 258.2300 ;
        RECT 984.6500 256.2300 986.6500 258.2300 ;
        RECT 1009.1000 249.1350 1011.1000 251.1350 ;
        RECT 1000.9500 249.1350 1002.9500 251.1350 ;
        RECT 992.8000 249.1350 994.8000 251.1350 ;
        RECT 984.6500 249.1350 986.6500 251.1350 ;
        RECT 992.8000 263.3250 994.8000 265.3250 ;
        RECT 984.6500 263.3250 986.6500 265.3250 ;
        RECT 1000.9500 263.3250 1002.9500 265.3250 ;
        RECT 1009.1000 263.3250 1011.1000 265.3250 ;
        RECT 984.6500 270.4200 986.6500 272.4200 ;
        RECT 992.8000 270.4200 994.8000 272.4200 ;
        RECT 1000.9500 270.4200 1002.9500 272.4200 ;
        RECT 1009.1000 270.4200 1011.1000 272.4200 ;
        RECT 984.6500 277.5150 986.6500 279.5150 ;
        RECT 992.8000 277.5150 994.8000 279.5150 ;
        RECT 1000.9500 277.5150 1002.9500 279.5150 ;
        RECT 1009.1000 277.5150 1011.1000 279.5150 ;
        RECT 1041.7000 256.2300 1043.7000 258.2300 ;
        RECT 1033.5500 256.2300 1035.5500 258.2300 ;
        RECT 1025.4000 256.2300 1027.4000 258.2300 ;
        RECT 1017.2500 256.2300 1019.2500 258.2300 ;
        RECT 1041.7000 249.1350 1043.7000 251.1350 ;
        RECT 1033.5500 249.1350 1035.5500 251.1350 ;
        RECT 1025.4000 249.1350 1027.4000 251.1350 ;
        RECT 1017.2500 249.1350 1019.2500 251.1350 ;
        RECT 1025.4000 263.3250 1027.4000 265.3250 ;
        RECT 1017.2500 263.3250 1019.2500 265.3250 ;
        RECT 1033.5500 263.3250 1035.5500 265.3250 ;
        RECT 1041.7000 263.3250 1043.7000 265.3250 ;
        RECT 1017.2500 270.4200 1019.2500 272.4200 ;
        RECT 1025.4000 270.4200 1027.4000 272.4200 ;
        RECT 1033.5500 270.4200 1035.5500 272.4200 ;
        RECT 1041.7000 270.4200 1043.7000 272.4200 ;
        RECT 1017.2500 277.5150 1019.2500 279.5150 ;
        RECT 1025.4000 277.5150 1027.4000 279.5150 ;
        RECT 1033.5500 277.5150 1035.5500 279.5150 ;
        RECT 1041.7000 277.5150 1043.7000 279.5150 ;
        RECT 1058.0000 220.7550 1060.0000 222.7550 ;
        RECT 1058.0000 213.6600 1060.0000 215.6600 ;
        RECT 1074.0000 220.7550 1076.0000 222.7550 ;
        RECT 1074.0000 213.6600 1076.0000 215.6600 ;
        RECT 1058.0000 227.8500 1060.0000 229.8500 ;
        RECT 1058.0000 234.9450 1060.0000 236.9450 ;
        RECT 1058.0000 242.0400 1060.0000 244.0400 ;
        RECT 1074.0000 234.9450 1076.0000 236.9450 ;
        RECT 1074.0000 227.8500 1076.0000 229.8500 ;
        RECT 1074.0000 242.0400 1076.0000 244.0400 ;
        RECT 1112.0000 213.6600 1114.0000 215.6600 ;
        RECT 1112.0000 220.7550 1114.0000 222.7550 ;
        RECT 1112.0000 234.9450 1114.0000 236.9450 ;
        RECT 1112.0000 227.8500 1114.0000 229.8500 ;
        RECT 1112.0000 242.0400 1114.0000 244.0400 ;
        RECT 1058.0000 256.2300 1060.0000 258.2300 ;
        RECT 1058.0000 249.1350 1060.0000 251.1350 ;
        RECT 1074.0000 249.1350 1076.0000 251.1350 ;
        RECT 1074.0000 256.2300 1076.0000 258.2300 ;
        RECT 1058.0000 270.4200 1060.0000 272.4200 ;
        RECT 1058.0000 263.3250 1060.0000 265.3250 ;
        RECT 1058.0000 277.5150 1060.0000 279.5150 ;
        RECT 1074.0000 270.4200 1076.0000 272.4200 ;
        RECT 1074.0000 263.3250 1076.0000 265.3250 ;
        RECT 1074.0000 277.5150 1076.0000 279.5150 ;
        RECT 1112.0000 249.1350 1114.0000 251.1350 ;
        RECT 1112.0000 256.2300 1114.0000 258.2300 ;
        RECT 1112.0000 270.4200 1114.0000 272.4200 ;
        RECT 1112.0000 263.3250 1114.0000 265.3250 ;
        RECT 1112.0000 277.5150 1114.0000 279.5150 ;
        RECT 699.4000 419.4150 701.4000 421.4150 ;
        RECT 626.0500 419.4150 628.0500 421.4150 ;
        RECT 617.9000 419.4150 619.9000 421.4150 ;
        RECT 609.7500 419.4150 611.7500 421.4150 ;
        RECT 601.6000 419.4150 603.6000 421.4150 ;
        RECT 593.4500 419.4150 595.4500 421.4150 ;
        RECT 585.3000 419.4150 587.3000 421.4150 ;
        RECT 577.1500 419.4150 579.1500 421.4150 ;
        RECT 569.0000 419.4150 571.0000 421.4150 ;
        RECT 560.8500 419.4150 562.8500 421.4150 ;
        RECT 658.6500 419.4150 660.6500 421.4150 ;
        RECT 650.5000 419.4150 652.5000 421.4150 ;
        RECT 642.3500 419.4150 644.3500 421.4150 ;
        RECT 634.2000 419.4150 636.2000 421.4150 ;
        RECT 666.8000 419.4150 668.8000 421.4150 ;
        RECT 674.9500 419.4150 676.9500 421.4150 ;
        RECT 683.1000 419.4150 685.1000 421.4150 ;
        RECT 691.2500 419.4150 693.2500 421.4150 ;
        RECT 764.6000 419.4150 766.6000 421.4150 ;
        RECT 756.4500 419.4150 758.4500 421.4150 ;
        RECT 748.3000 419.4150 750.3000 421.4150 ;
        RECT 740.1500 419.4150 742.1500 421.4150 ;
        RECT 732.0000 419.4150 734.0000 421.4150 ;
        RECT 723.8500 419.4150 725.8500 421.4150 ;
        RECT 715.7000 419.4150 717.7000 421.4150 ;
        RECT 707.5500 419.4150 709.5500 421.4150 ;
        RECT 805.3500 419.4150 807.3500 421.4150 ;
        RECT 797.2000 419.4150 799.2000 421.4150 ;
        RECT 789.0500 419.4150 791.0500 421.4150 ;
        RECT 780.9000 419.4150 782.9000 421.4150 ;
        RECT 772.7500 419.4150 774.7500 421.4150 ;
        RECT 813.5000 419.4150 815.5000 421.4150 ;
        RECT 821.6500 419.4150 823.6500 421.4150 ;
        RECT 829.8000 419.4150 831.8000 421.4150 ;
        RECT 837.9500 419.4150 839.9500 421.4150 ;
        RECT 699.4000 348.4650 701.4000 350.4650 ;
        RECT 699.4000 341.3700 701.4000 343.3700 ;
        RECT 699.4000 334.2750 701.4000 336.2750 ;
        RECT 699.4000 327.1800 701.4000 329.1800 ;
        RECT 699.4000 320.0850 701.4000 322.0850 ;
        RECT 699.4000 312.9900 701.4000 314.9900 ;
        RECT 699.4000 305.8950 701.4000 307.8950 ;
        RECT 699.4000 298.8000 701.4000 300.8000 ;
        RECT 699.4000 291.7050 701.4000 293.7050 ;
        RECT 699.4000 284.6100 701.4000 286.6100 ;
        RECT 699.4000 355.5600 701.4000 357.5600 ;
        RECT 699.4000 362.6550 701.4000 364.6550 ;
        RECT 699.4000 369.7500 701.4000 371.7500 ;
        RECT 699.4000 376.8450 701.4000 378.8450 ;
        RECT 699.4000 383.9400 701.4000 385.9400 ;
        RECT 699.4000 391.0350 701.4000 393.0350 ;
        RECT 699.4000 398.1300 701.4000 400.1300 ;
        RECT 699.4000 405.2250 701.4000 407.2250 ;
        RECT 699.4000 412.3200 701.4000 414.3200 ;
        RECT 626.0500 348.4650 628.0500 350.4650 ;
        RECT 617.9000 348.4650 619.9000 350.4650 ;
        RECT 609.7500 348.4650 611.7500 350.4650 ;
        RECT 601.6000 348.4650 603.6000 350.4650 ;
        RECT 593.4500 348.4650 595.4500 350.4650 ;
        RECT 585.3000 348.4650 587.3000 350.4650 ;
        RECT 577.1500 348.4650 579.1500 350.4650 ;
        RECT 569.0000 348.4650 571.0000 350.4650 ;
        RECT 560.8500 348.4650 562.8500 350.4650 ;
        RECT 658.6500 348.4650 660.6500 350.4650 ;
        RECT 650.5000 348.4650 652.5000 350.4650 ;
        RECT 642.3500 348.4650 644.3500 350.4650 ;
        RECT 634.2000 348.4650 636.2000 350.4650 ;
        RECT 666.8000 348.4650 668.8000 350.4650 ;
        RECT 674.9500 348.4650 676.9500 350.4650 ;
        RECT 683.1000 348.4650 685.1000 350.4650 ;
        RECT 691.2500 348.4650 693.2500 350.4650 ;
        RECT 593.4500 284.6100 595.4500 286.6100 ;
        RECT 593.4500 291.7050 595.4500 293.7050 ;
        RECT 593.4500 298.8000 595.4500 300.8000 ;
        RECT 593.4500 305.8950 595.4500 307.8950 ;
        RECT 593.4500 312.9900 595.4500 314.9900 ;
        RECT 585.3000 291.7050 587.3000 293.7050 ;
        RECT 577.1500 291.7050 579.1500 293.7050 ;
        RECT 569.0000 291.7050 571.0000 293.7050 ;
        RECT 560.8500 291.7050 562.8500 293.7050 ;
        RECT 585.3000 284.6100 587.3000 286.6100 ;
        RECT 577.1500 284.6100 579.1500 286.6100 ;
        RECT 569.0000 284.6100 571.0000 286.6100 ;
        RECT 560.8500 284.6100 562.8500 286.6100 ;
        RECT 569.0000 298.8000 571.0000 300.8000 ;
        RECT 560.8500 298.8000 562.8500 300.8000 ;
        RECT 577.1500 298.8000 579.1500 300.8000 ;
        RECT 585.3000 298.8000 587.3000 300.8000 ;
        RECT 560.8500 305.8950 562.8500 307.8950 ;
        RECT 569.0000 305.8950 571.0000 307.8950 ;
        RECT 577.1500 305.8950 579.1500 307.8950 ;
        RECT 585.3000 305.8950 587.3000 307.8950 ;
        RECT 560.8500 312.9900 562.8500 314.9900 ;
        RECT 569.0000 312.9900 571.0000 314.9900 ;
        RECT 577.1500 312.9900 579.1500 314.9900 ;
        RECT 585.3000 312.9900 587.3000 314.9900 ;
        RECT 626.0500 291.7050 628.0500 293.7050 ;
        RECT 617.9000 291.7050 619.9000 293.7050 ;
        RECT 609.7500 291.7050 611.7500 293.7050 ;
        RECT 601.6000 291.7050 603.6000 293.7050 ;
        RECT 626.0500 284.6100 628.0500 286.6100 ;
        RECT 617.9000 284.6100 619.9000 286.6100 ;
        RECT 609.7500 284.6100 611.7500 286.6100 ;
        RECT 601.6000 284.6100 603.6000 286.6100 ;
        RECT 609.7500 298.8000 611.7500 300.8000 ;
        RECT 601.6000 298.8000 603.6000 300.8000 ;
        RECT 617.9000 298.8000 619.9000 300.8000 ;
        RECT 626.0500 298.8000 628.0500 300.8000 ;
        RECT 601.6000 305.8950 603.6000 307.8950 ;
        RECT 609.7500 305.8950 611.7500 307.8950 ;
        RECT 617.9000 305.8950 619.9000 307.8950 ;
        RECT 626.0500 305.8950 628.0500 307.8950 ;
        RECT 601.6000 312.9900 603.6000 314.9900 ;
        RECT 609.7500 312.9900 611.7500 314.9900 ;
        RECT 617.9000 312.9900 619.9000 314.9900 ;
        RECT 626.0500 312.9900 628.0500 314.9900 ;
        RECT 593.4500 320.0850 595.4500 322.0850 ;
        RECT 593.4500 327.1800 595.4500 329.1800 ;
        RECT 593.4500 334.2750 595.4500 336.2750 ;
        RECT 593.4500 341.3700 595.4500 343.3700 ;
        RECT 585.3000 327.1800 587.3000 329.1800 ;
        RECT 577.1500 327.1800 579.1500 329.1800 ;
        RECT 569.0000 327.1800 571.0000 329.1800 ;
        RECT 560.8500 327.1800 562.8500 329.1800 ;
        RECT 585.3000 320.0850 587.3000 322.0850 ;
        RECT 577.1500 320.0850 579.1500 322.0850 ;
        RECT 569.0000 320.0850 571.0000 322.0850 ;
        RECT 560.8500 320.0850 562.8500 322.0850 ;
        RECT 569.0000 341.3700 571.0000 343.3700 ;
        RECT 560.8500 341.3700 562.8500 343.3700 ;
        RECT 585.3000 334.2750 587.3000 336.2750 ;
        RECT 577.1500 334.2750 579.1500 336.2750 ;
        RECT 569.0000 334.2750 571.0000 336.2750 ;
        RECT 560.8500 334.2750 562.8500 336.2750 ;
        RECT 577.1500 341.3700 579.1500 343.3700 ;
        RECT 585.3000 341.3700 587.3000 343.3700 ;
        RECT 626.0500 327.1800 628.0500 329.1800 ;
        RECT 617.9000 327.1800 619.9000 329.1800 ;
        RECT 609.7500 327.1800 611.7500 329.1800 ;
        RECT 601.6000 327.1800 603.6000 329.1800 ;
        RECT 626.0500 320.0850 628.0500 322.0850 ;
        RECT 617.9000 320.0850 619.9000 322.0850 ;
        RECT 609.7500 320.0850 611.7500 322.0850 ;
        RECT 601.6000 320.0850 603.6000 322.0850 ;
        RECT 609.7500 341.3700 611.7500 343.3700 ;
        RECT 601.6000 341.3700 603.6000 343.3700 ;
        RECT 626.0500 334.2750 628.0500 336.2750 ;
        RECT 617.9000 334.2750 619.9000 336.2750 ;
        RECT 609.7500 334.2750 611.7500 336.2750 ;
        RECT 601.6000 334.2750 603.6000 336.2750 ;
        RECT 617.9000 341.3700 619.9000 343.3700 ;
        RECT 626.0500 341.3700 628.0500 343.3700 ;
        RECT 658.6500 291.7050 660.6500 293.7050 ;
        RECT 650.5000 291.7050 652.5000 293.7050 ;
        RECT 642.3500 291.7050 644.3500 293.7050 ;
        RECT 634.2000 291.7050 636.2000 293.7050 ;
        RECT 658.6500 284.6100 660.6500 286.6100 ;
        RECT 650.5000 284.6100 652.5000 286.6100 ;
        RECT 642.3500 284.6100 644.3500 286.6100 ;
        RECT 634.2000 284.6100 636.2000 286.6100 ;
        RECT 642.3500 298.8000 644.3500 300.8000 ;
        RECT 634.2000 298.8000 636.2000 300.8000 ;
        RECT 650.5000 298.8000 652.5000 300.8000 ;
        RECT 658.6500 298.8000 660.6500 300.8000 ;
        RECT 634.2000 305.8950 636.2000 307.8950 ;
        RECT 642.3500 305.8950 644.3500 307.8950 ;
        RECT 650.5000 305.8950 652.5000 307.8950 ;
        RECT 658.6500 305.8950 660.6500 307.8950 ;
        RECT 634.2000 312.9900 636.2000 314.9900 ;
        RECT 642.3500 312.9900 644.3500 314.9900 ;
        RECT 650.5000 312.9900 652.5000 314.9900 ;
        RECT 658.6500 312.9900 660.6500 314.9900 ;
        RECT 691.2500 291.7050 693.2500 293.7050 ;
        RECT 683.1000 291.7050 685.1000 293.7050 ;
        RECT 674.9500 291.7050 676.9500 293.7050 ;
        RECT 666.8000 291.7050 668.8000 293.7050 ;
        RECT 691.2500 284.6100 693.2500 286.6100 ;
        RECT 683.1000 284.6100 685.1000 286.6100 ;
        RECT 674.9500 284.6100 676.9500 286.6100 ;
        RECT 666.8000 284.6100 668.8000 286.6100 ;
        RECT 674.9500 298.8000 676.9500 300.8000 ;
        RECT 666.8000 298.8000 668.8000 300.8000 ;
        RECT 683.1000 298.8000 685.1000 300.8000 ;
        RECT 691.2500 298.8000 693.2500 300.8000 ;
        RECT 666.8000 305.8950 668.8000 307.8950 ;
        RECT 674.9500 305.8950 676.9500 307.8950 ;
        RECT 683.1000 305.8950 685.1000 307.8950 ;
        RECT 691.2500 305.8950 693.2500 307.8950 ;
        RECT 666.8000 312.9900 668.8000 314.9900 ;
        RECT 674.9500 312.9900 676.9500 314.9900 ;
        RECT 683.1000 312.9900 685.1000 314.9900 ;
        RECT 691.2500 312.9900 693.2500 314.9900 ;
        RECT 658.6500 327.1800 660.6500 329.1800 ;
        RECT 650.5000 327.1800 652.5000 329.1800 ;
        RECT 642.3500 327.1800 644.3500 329.1800 ;
        RECT 634.2000 327.1800 636.2000 329.1800 ;
        RECT 658.6500 320.0850 660.6500 322.0850 ;
        RECT 650.5000 320.0850 652.5000 322.0850 ;
        RECT 642.3500 320.0850 644.3500 322.0850 ;
        RECT 634.2000 320.0850 636.2000 322.0850 ;
        RECT 642.3500 341.3700 644.3500 343.3700 ;
        RECT 634.2000 341.3700 636.2000 343.3700 ;
        RECT 658.6500 334.2750 660.6500 336.2750 ;
        RECT 650.5000 334.2750 652.5000 336.2750 ;
        RECT 642.3500 334.2750 644.3500 336.2750 ;
        RECT 634.2000 334.2750 636.2000 336.2750 ;
        RECT 650.5000 341.3700 652.5000 343.3700 ;
        RECT 658.6500 341.3700 660.6500 343.3700 ;
        RECT 691.2500 327.1800 693.2500 329.1800 ;
        RECT 683.1000 327.1800 685.1000 329.1800 ;
        RECT 674.9500 327.1800 676.9500 329.1800 ;
        RECT 666.8000 327.1800 668.8000 329.1800 ;
        RECT 691.2500 320.0850 693.2500 322.0850 ;
        RECT 683.1000 320.0850 685.1000 322.0850 ;
        RECT 674.9500 320.0850 676.9500 322.0850 ;
        RECT 666.8000 320.0850 668.8000 322.0850 ;
        RECT 674.9500 341.3700 676.9500 343.3700 ;
        RECT 666.8000 341.3700 668.8000 343.3700 ;
        RECT 691.2500 334.2750 693.2500 336.2750 ;
        RECT 683.1000 334.2750 685.1000 336.2750 ;
        RECT 674.9500 334.2750 676.9500 336.2750 ;
        RECT 666.8000 334.2750 668.8000 336.2750 ;
        RECT 683.1000 341.3700 685.1000 343.3700 ;
        RECT 691.2500 341.3700 693.2500 343.3700 ;
        RECT 560.8500 383.9400 562.8500 385.9400 ;
        RECT 569.0000 383.9400 571.0000 385.9400 ;
        RECT 577.1500 383.9400 579.1500 385.9400 ;
        RECT 585.3000 383.9400 587.3000 385.9400 ;
        RECT 593.4500 383.9400 595.4500 385.9400 ;
        RECT 601.6000 383.9400 603.6000 385.9400 ;
        RECT 609.7500 383.9400 611.7500 385.9400 ;
        RECT 617.9000 383.9400 619.9000 385.9400 ;
        RECT 626.0500 383.9400 628.0500 385.9400 ;
        RECT 593.4500 355.5600 595.4500 357.5600 ;
        RECT 593.4500 362.6550 595.4500 364.6550 ;
        RECT 593.4500 369.7500 595.4500 371.7500 ;
        RECT 593.4500 376.8450 595.4500 378.8450 ;
        RECT 585.3000 362.6550 587.3000 364.6550 ;
        RECT 577.1500 362.6550 579.1500 364.6550 ;
        RECT 569.0000 362.6550 571.0000 364.6550 ;
        RECT 560.8500 362.6550 562.8500 364.6550 ;
        RECT 585.3000 355.5600 587.3000 357.5600 ;
        RECT 577.1500 355.5600 579.1500 357.5600 ;
        RECT 569.0000 355.5600 571.0000 357.5600 ;
        RECT 560.8500 355.5600 562.8500 357.5600 ;
        RECT 569.0000 376.8450 571.0000 378.8450 ;
        RECT 560.8500 376.8450 562.8500 378.8450 ;
        RECT 585.3000 369.7500 587.3000 371.7500 ;
        RECT 577.1500 369.7500 579.1500 371.7500 ;
        RECT 569.0000 369.7500 571.0000 371.7500 ;
        RECT 560.8500 369.7500 562.8500 371.7500 ;
        RECT 577.1500 376.8450 579.1500 378.8450 ;
        RECT 585.3000 376.8450 587.3000 378.8450 ;
        RECT 626.0500 362.6550 628.0500 364.6550 ;
        RECT 617.9000 362.6550 619.9000 364.6550 ;
        RECT 609.7500 362.6550 611.7500 364.6550 ;
        RECT 601.6000 362.6550 603.6000 364.6550 ;
        RECT 626.0500 355.5600 628.0500 357.5600 ;
        RECT 617.9000 355.5600 619.9000 357.5600 ;
        RECT 609.7500 355.5600 611.7500 357.5600 ;
        RECT 601.6000 355.5600 603.6000 357.5600 ;
        RECT 609.7500 376.8450 611.7500 378.8450 ;
        RECT 601.6000 376.8450 603.6000 378.8450 ;
        RECT 626.0500 369.7500 628.0500 371.7500 ;
        RECT 617.9000 369.7500 619.9000 371.7500 ;
        RECT 609.7500 369.7500 611.7500 371.7500 ;
        RECT 601.6000 369.7500 603.6000 371.7500 ;
        RECT 617.9000 376.8450 619.9000 378.8450 ;
        RECT 626.0500 376.8450 628.0500 378.8450 ;
        RECT 593.4500 391.0350 595.4500 393.0350 ;
        RECT 593.4500 398.1300 595.4500 400.1300 ;
        RECT 593.4500 405.2250 595.4500 407.2250 ;
        RECT 593.4500 412.3200 595.4500 414.3200 ;
        RECT 585.3000 398.1300 587.3000 400.1300 ;
        RECT 577.1500 398.1300 579.1500 400.1300 ;
        RECT 569.0000 398.1300 571.0000 400.1300 ;
        RECT 560.8500 398.1300 562.8500 400.1300 ;
        RECT 585.3000 391.0350 587.3000 393.0350 ;
        RECT 577.1500 391.0350 579.1500 393.0350 ;
        RECT 569.0000 391.0350 571.0000 393.0350 ;
        RECT 560.8500 391.0350 562.8500 393.0350 ;
        RECT 569.0000 412.3200 571.0000 414.3200 ;
        RECT 560.8500 412.3200 562.8500 414.3200 ;
        RECT 585.3000 405.2250 587.3000 407.2250 ;
        RECT 577.1500 405.2250 579.1500 407.2250 ;
        RECT 569.0000 405.2250 571.0000 407.2250 ;
        RECT 560.8500 405.2250 562.8500 407.2250 ;
        RECT 577.1500 412.3200 579.1500 414.3200 ;
        RECT 585.3000 412.3200 587.3000 414.3200 ;
        RECT 626.0500 398.1300 628.0500 400.1300 ;
        RECT 617.9000 398.1300 619.9000 400.1300 ;
        RECT 609.7500 398.1300 611.7500 400.1300 ;
        RECT 601.6000 398.1300 603.6000 400.1300 ;
        RECT 626.0500 391.0350 628.0500 393.0350 ;
        RECT 617.9000 391.0350 619.9000 393.0350 ;
        RECT 609.7500 391.0350 611.7500 393.0350 ;
        RECT 601.6000 391.0350 603.6000 393.0350 ;
        RECT 609.7500 412.3200 611.7500 414.3200 ;
        RECT 601.6000 412.3200 603.6000 414.3200 ;
        RECT 626.0500 405.2250 628.0500 407.2250 ;
        RECT 617.9000 405.2250 619.9000 407.2250 ;
        RECT 609.7500 405.2250 611.7500 407.2250 ;
        RECT 601.6000 405.2250 603.6000 407.2250 ;
        RECT 617.9000 412.3200 619.9000 414.3200 ;
        RECT 626.0500 412.3200 628.0500 414.3200 ;
        RECT 634.2000 383.9400 636.2000 385.9400 ;
        RECT 642.3500 383.9400 644.3500 385.9400 ;
        RECT 650.5000 383.9400 652.5000 385.9400 ;
        RECT 658.6500 383.9400 660.6500 385.9400 ;
        RECT 666.8000 383.9400 668.8000 385.9400 ;
        RECT 674.9500 383.9400 676.9500 385.9400 ;
        RECT 683.1000 383.9400 685.1000 385.9400 ;
        RECT 691.2500 383.9400 693.2500 385.9400 ;
        RECT 658.6500 362.6550 660.6500 364.6550 ;
        RECT 650.5000 362.6550 652.5000 364.6550 ;
        RECT 642.3500 362.6550 644.3500 364.6550 ;
        RECT 634.2000 362.6550 636.2000 364.6550 ;
        RECT 658.6500 355.5600 660.6500 357.5600 ;
        RECT 650.5000 355.5600 652.5000 357.5600 ;
        RECT 642.3500 355.5600 644.3500 357.5600 ;
        RECT 634.2000 355.5600 636.2000 357.5600 ;
        RECT 642.3500 376.8450 644.3500 378.8450 ;
        RECT 634.2000 376.8450 636.2000 378.8450 ;
        RECT 658.6500 369.7500 660.6500 371.7500 ;
        RECT 650.5000 369.7500 652.5000 371.7500 ;
        RECT 642.3500 369.7500 644.3500 371.7500 ;
        RECT 634.2000 369.7500 636.2000 371.7500 ;
        RECT 650.5000 376.8450 652.5000 378.8450 ;
        RECT 658.6500 376.8450 660.6500 378.8450 ;
        RECT 691.2500 362.6550 693.2500 364.6550 ;
        RECT 683.1000 362.6550 685.1000 364.6550 ;
        RECT 674.9500 362.6550 676.9500 364.6550 ;
        RECT 666.8000 362.6550 668.8000 364.6550 ;
        RECT 691.2500 355.5600 693.2500 357.5600 ;
        RECT 683.1000 355.5600 685.1000 357.5600 ;
        RECT 674.9500 355.5600 676.9500 357.5600 ;
        RECT 666.8000 355.5600 668.8000 357.5600 ;
        RECT 674.9500 376.8450 676.9500 378.8450 ;
        RECT 666.8000 376.8450 668.8000 378.8450 ;
        RECT 691.2500 369.7500 693.2500 371.7500 ;
        RECT 683.1000 369.7500 685.1000 371.7500 ;
        RECT 674.9500 369.7500 676.9500 371.7500 ;
        RECT 666.8000 369.7500 668.8000 371.7500 ;
        RECT 683.1000 376.8450 685.1000 378.8450 ;
        RECT 691.2500 376.8450 693.2500 378.8450 ;
        RECT 658.6500 398.1300 660.6500 400.1300 ;
        RECT 650.5000 398.1300 652.5000 400.1300 ;
        RECT 642.3500 398.1300 644.3500 400.1300 ;
        RECT 634.2000 398.1300 636.2000 400.1300 ;
        RECT 658.6500 391.0350 660.6500 393.0350 ;
        RECT 650.5000 391.0350 652.5000 393.0350 ;
        RECT 642.3500 391.0350 644.3500 393.0350 ;
        RECT 634.2000 391.0350 636.2000 393.0350 ;
        RECT 642.3500 412.3200 644.3500 414.3200 ;
        RECT 634.2000 412.3200 636.2000 414.3200 ;
        RECT 658.6500 405.2250 660.6500 407.2250 ;
        RECT 650.5000 405.2250 652.5000 407.2250 ;
        RECT 642.3500 405.2250 644.3500 407.2250 ;
        RECT 634.2000 405.2250 636.2000 407.2250 ;
        RECT 650.5000 412.3200 652.5000 414.3200 ;
        RECT 658.6500 412.3200 660.6500 414.3200 ;
        RECT 691.2500 398.1300 693.2500 400.1300 ;
        RECT 683.1000 398.1300 685.1000 400.1300 ;
        RECT 674.9500 398.1300 676.9500 400.1300 ;
        RECT 666.8000 398.1300 668.8000 400.1300 ;
        RECT 691.2500 391.0350 693.2500 393.0350 ;
        RECT 683.1000 391.0350 685.1000 393.0350 ;
        RECT 674.9500 391.0350 676.9500 393.0350 ;
        RECT 666.8000 391.0350 668.8000 393.0350 ;
        RECT 674.9500 412.3200 676.9500 414.3200 ;
        RECT 666.8000 412.3200 668.8000 414.3200 ;
        RECT 691.2500 405.2250 693.2500 407.2250 ;
        RECT 683.1000 405.2250 685.1000 407.2250 ;
        RECT 674.9500 405.2250 676.9500 407.2250 ;
        RECT 666.8000 405.2250 668.8000 407.2250 ;
        RECT 683.1000 412.3200 685.1000 414.3200 ;
        RECT 691.2500 412.3200 693.2500 414.3200 ;
        RECT 764.6000 348.4650 766.6000 350.4650 ;
        RECT 756.4500 348.4650 758.4500 350.4650 ;
        RECT 748.3000 348.4650 750.3000 350.4650 ;
        RECT 740.1500 348.4650 742.1500 350.4650 ;
        RECT 732.0000 348.4650 734.0000 350.4650 ;
        RECT 723.8500 348.4650 725.8500 350.4650 ;
        RECT 715.7000 348.4650 717.7000 350.4650 ;
        RECT 707.5500 348.4650 709.5500 350.4650 ;
        RECT 805.3500 348.4650 807.3500 350.4650 ;
        RECT 797.2000 348.4650 799.2000 350.4650 ;
        RECT 789.0500 348.4650 791.0500 350.4650 ;
        RECT 780.9000 348.4650 782.9000 350.4650 ;
        RECT 772.7500 348.4650 774.7500 350.4650 ;
        RECT 813.5000 348.4650 815.5000 350.4650 ;
        RECT 821.6500 348.4650 823.6500 350.4650 ;
        RECT 829.8000 348.4650 831.8000 350.4650 ;
        RECT 837.9500 348.4650 839.9500 350.4650 ;
        RECT 732.0000 291.7050 734.0000 293.7050 ;
        RECT 723.8500 291.7050 725.8500 293.7050 ;
        RECT 715.7000 291.7050 717.7000 293.7050 ;
        RECT 707.5500 291.7050 709.5500 293.7050 ;
        RECT 732.0000 284.6100 734.0000 286.6100 ;
        RECT 723.8500 284.6100 725.8500 286.6100 ;
        RECT 715.7000 284.6100 717.7000 286.6100 ;
        RECT 707.5500 284.6100 709.5500 286.6100 ;
        RECT 715.7000 298.8000 717.7000 300.8000 ;
        RECT 707.5500 298.8000 709.5500 300.8000 ;
        RECT 723.8500 298.8000 725.8500 300.8000 ;
        RECT 732.0000 298.8000 734.0000 300.8000 ;
        RECT 707.5500 305.8950 709.5500 307.8950 ;
        RECT 715.7000 305.8950 717.7000 307.8950 ;
        RECT 723.8500 305.8950 725.8500 307.8950 ;
        RECT 732.0000 305.8950 734.0000 307.8950 ;
        RECT 707.5500 312.9900 709.5500 314.9900 ;
        RECT 715.7000 312.9900 717.7000 314.9900 ;
        RECT 723.8500 312.9900 725.8500 314.9900 ;
        RECT 732.0000 312.9900 734.0000 314.9900 ;
        RECT 764.6000 291.7050 766.6000 293.7050 ;
        RECT 756.4500 291.7050 758.4500 293.7050 ;
        RECT 748.3000 291.7050 750.3000 293.7050 ;
        RECT 740.1500 291.7050 742.1500 293.7050 ;
        RECT 764.6000 284.6100 766.6000 286.6100 ;
        RECT 756.4500 284.6100 758.4500 286.6100 ;
        RECT 748.3000 284.6100 750.3000 286.6100 ;
        RECT 740.1500 284.6100 742.1500 286.6100 ;
        RECT 748.3000 298.8000 750.3000 300.8000 ;
        RECT 740.1500 298.8000 742.1500 300.8000 ;
        RECT 756.4500 298.8000 758.4500 300.8000 ;
        RECT 764.6000 298.8000 766.6000 300.8000 ;
        RECT 740.1500 305.8950 742.1500 307.8950 ;
        RECT 748.3000 305.8950 750.3000 307.8950 ;
        RECT 756.4500 305.8950 758.4500 307.8950 ;
        RECT 764.6000 305.8950 766.6000 307.8950 ;
        RECT 740.1500 312.9900 742.1500 314.9900 ;
        RECT 748.3000 312.9900 750.3000 314.9900 ;
        RECT 756.4500 312.9900 758.4500 314.9900 ;
        RECT 764.6000 312.9900 766.6000 314.9900 ;
        RECT 732.0000 327.1800 734.0000 329.1800 ;
        RECT 723.8500 327.1800 725.8500 329.1800 ;
        RECT 715.7000 327.1800 717.7000 329.1800 ;
        RECT 707.5500 327.1800 709.5500 329.1800 ;
        RECT 732.0000 320.0850 734.0000 322.0850 ;
        RECT 723.8500 320.0850 725.8500 322.0850 ;
        RECT 715.7000 320.0850 717.7000 322.0850 ;
        RECT 707.5500 320.0850 709.5500 322.0850 ;
        RECT 715.7000 341.3700 717.7000 343.3700 ;
        RECT 707.5500 341.3700 709.5500 343.3700 ;
        RECT 732.0000 334.2750 734.0000 336.2750 ;
        RECT 723.8500 334.2750 725.8500 336.2750 ;
        RECT 715.7000 334.2750 717.7000 336.2750 ;
        RECT 707.5500 334.2750 709.5500 336.2750 ;
        RECT 723.8500 341.3700 725.8500 343.3700 ;
        RECT 732.0000 341.3700 734.0000 343.3700 ;
        RECT 764.6000 327.1800 766.6000 329.1800 ;
        RECT 756.4500 327.1800 758.4500 329.1800 ;
        RECT 748.3000 327.1800 750.3000 329.1800 ;
        RECT 740.1500 327.1800 742.1500 329.1800 ;
        RECT 764.6000 320.0850 766.6000 322.0850 ;
        RECT 756.4500 320.0850 758.4500 322.0850 ;
        RECT 748.3000 320.0850 750.3000 322.0850 ;
        RECT 740.1500 320.0850 742.1500 322.0850 ;
        RECT 748.3000 341.3700 750.3000 343.3700 ;
        RECT 740.1500 341.3700 742.1500 343.3700 ;
        RECT 764.6000 334.2750 766.6000 336.2750 ;
        RECT 756.4500 334.2750 758.4500 336.2750 ;
        RECT 748.3000 334.2750 750.3000 336.2750 ;
        RECT 740.1500 334.2750 742.1500 336.2750 ;
        RECT 756.4500 341.3700 758.4500 343.3700 ;
        RECT 764.6000 341.3700 766.6000 343.3700 ;
        RECT 797.2000 291.7050 799.2000 293.7050 ;
        RECT 789.0500 291.7050 791.0500 293.7050 ;
        RECT 780.9000 291.7050 782.9000 293.7050 ;
        RECT 772.7500 291.7050 774.7500 293.7050 ;
        RECT 797.2000 284.6100 799.2000 286.6100 ;
        RECT 789.0500 284.6100 791.0500 286.6100 ;
        RECT 780.9000 284.6100 782.9000 286.6100 ;
        RECT 772.7500 284.6100 774.7500 286.6100 ;
        RECT 780.9000 298.8000 782.9000 300.8000 ;
        RECT 772.7500 298.8000 774.7500 300.8000 ;
        RECT 789.0500 298.8000 791.0500 300.8000 ;
        RECT 797.2000 298.8000 799.2000 300.8000 ;
        RECT 772.7500 305.8950 774.7500 307.8950 ;
        RECT 780.9000 305.8950 782.9000 307.8950 ;
        RECT 789.0500 305.8950 791.0500 307.8950 ;
        RECT 797.2000 305.8950 799.2000 307.8950 ;
        RECT 772.7500 312.9900 774.7500 314.9900 ;
        RECT 780.9000 312.9900 782.9000 314.9900 ;
        RECT 789.0500 312.9900 791.0500 314.9900 ;
        RECT 797.2000 312.9900 799.2000 314.9900 ;
        RECT 837.9500 284.6100 839.9500 286.6100 ;
        RECT 829.8000 284.6100 831.8000 286.6100 ;
        RECT 821.6500 284.6100 823.6500 286.6100 ;
        RECT 813.5000 284.6100 815.5000 286.6100 ;
        RECT 805.3500 284.6100 807.3500 286.6100 ;
        RECT 805.3500 291.7050 807.3500 293.7050 ;
        RECT 813.5000 291.7050 815.5000 293.7050 ;
        RECT 821.6500 291.7050 823.6500 293.7050 ;
        RECT 829.8000 291.7050 831.8000 293.7050 ;
        RECT 837.9500 291.7050 839.9500 293.7050 ;
        RECT 821.6500 298.8000 823.6500 300.8000 ;
        RECT 821.6500 305.8950 823.6500 307.8950 ;
        RECT 821.6500 312.9900 823.6500 314.9900 ;
        RECT 813.5000 312.9900 815.5000 314.9900 ;
        RECT 805.3500 312.9900 807.3500 314.9900 ;
        RECT 813.5000 305.8950 815.5000 307.8950 ;
        RECT 805.3500 305.8950 807.3500 307.8950 ;
        RECT 813.5000 298.8000 815.5000 300.8000 ;
        RECT 805.3500 298.8000 807.3500 300.8000 ;
        RECT 837.9500 312.9900 839.9500 314.9900 ;
        RECT 829.8000 312.9900 831.8000 314.9900 ;
        RECT 837.9500 305.8950 839.9500 307.8950 ;
        RECT 829.8000 305.8950 831.8000 307.8950 ;
        RECT 837.9500 298.8000 839.9500 300.8000 ;
        RECT 829.8000 298.8000 831.8000 300.8000 ;
        RECT 797.2000 327.1800 799.2000 329.1800 ;
        RECT 789.0500 327.1800 791.0500 329.1800 ;
        RECT 780.9000 327.1800 782.9000 329.1800 ;
        RECT 772.7500 327.1800 774.7500 329.1800 ;
        RECT 797.2000 320.0850 799.2000 322.0850 ;
        RECT 789.0500 320.0850 791.0500 322.0850 ;
        RECT 780.9000 320.0850 782.9000 322.0850 ;
        RECT 772.7500 320.0850 774.7500 322.0850 ;
        RECT 780.9000 341.3700 782.9000 343.3700 ;
        RECT 772.7500 341.3700 774.7500 343.3700 ;
        RECT 797.2000 334.2750 799.2000 336.2750 ;
        RECT 789.0500 334.2750 791.0500 336.2750 ;
        RECT 780.9000 334.2750 782.9000 336.2750 ;
        RECT 772.7500 334.2750 774.7500 336.2750 ;
        RECT 789.0500 341.3700 791.0500 343.3700 ;
        RECT 797.2000 341.3700 799.2000 343.3700 ;
        RECT 837.9500 327.1800 839.9500 329.1800 ;
        RECT 829.8000 327.1800 831.8000 329.1800 ;
        RECT 821.6500 327.1800 823.6500 329.1800 ;
        RECT 813.5000 327.1800 815.5000 329.1800 ;
        RECT 805.3500 327.1800 807.3500 329.1800 ;
        RECT 837.9500 320.0850 839.9500 322.0850 ;
        RECT 829.8000 320.0850 831.8000 322.0850 ;
        RECT 821.6500 320.0850 823.6500 322.0850 ;
        RECT 813.5000 320.0850 815.5000 322.0850 ;
        RECT 805.3500 320.0850 807.3500 322.0850 ;
        RECT 805.3500 334.2750 807.3500 336.2750 ;
        RECT 813.5000 334.2750 815.5000 336.2750 ;
        RECT 821.6500 334.2750 823.6500 336.2750 ;
        RECT 829.8000 334.2750 831.8000 336.2750 ;
        RECT 837.9500 334.2750 839.9500 336.2750 ;
        RECT 805.3500 341.3700 807.3500 343.3700 ;
        RECT 813.5000 341.3700 815.5000 343.3700 ;
        RECT 821.6500 341.3700 823.6500 343.3700 ;
        RECT 829.8000 341.3700 831.8000 343.3700 ;
        RECT 837.9500 341.3700 839.9500 343.3700 ;
        RECT 707.5500 383.9400 709.5500 385.9400 ;
        RECT 715.7000 383.9400 717.7000 385.9400 ;
        RECT 723.8500 383.9400 725.8500 385.9400 ;
        RECT 732.0000 383.9400 734.0000 385.9400 ;
        RECT 740.1500 383.9400 742.1500 385.9400 ;
        RECT 748.3000 383.9400 750.3000 385.9400 ;
        RECT 756.4500 383.9400 758.4500 385.9400 ;
        RECT 764.6000 383.9400 766.6000 385.9400 ;
        RECT 732.0000 362.6550 734.0000 364.6550 ;
        RECT 723.8500 362.6550 725.8500 364.6550 ;
        RECT 715.7000 362.6550 717.7000 364.6550 ;
        RECT 707.5500 362.6550 709.5500 364.6550 ;
        RECT 732.0000 355.5600 734.0000 357.5600 ;
        RECT 723.8500 355.5600 725.8500 357.5600 ;
        RECT 715.7000 355.5600 717.7000 357.5600 ;
        RECT 707.5500 355.5600 709.5500 357.5600 ;
        RECT 715.7000 376.8450 717.7000 378.8450 ;
        RECT 707.5500 376.8450 709.5500 378.8450 ;
        RECT 732.0000 369.7500 734.0000 371.7500 ;
        RECT 723.8500 369.7500 725.8500 371.7500 ;
        RECT 715.7000 369.7500 717.7000 371.7500 ;
        RECT 707.5500 369.7500 709.5500 371.7500 ;
        RECT 723.8500 376.8450 725.8500 378.8450 ;
        RECT 732.0000 376.8450 734.0000 378.8450 ;
        RECT 764.6000 362.6550 766.6000 364.6550 ;
        RECT 756.4500 362.6550 758.4500 364.6550 ;
        RECT 748.3000 362.6550 750.3000 364.6550 ;
        RECT 740.1500 362.6550 742.1500 364.6550 ;
        RECT 764.6000 355.5600 766.6000 357.5600 ;
        RECT 756.4500 355.5600 758.4500 357.5600 ;
        RECT 748.3000 355.5600 750.3000 357.5600 ;
        RECT 740.1500 355.5600 742.1500 357.5600 ;
        RECT 748.3000 376.8450 750.3000 378.8450 ;
        RECT 740.1500 376.8450 742.1500 378.8450 ;
        RECT 764.6000 369.7500 766.6000 371.7500 ;
        RECT 756.4500 369.7500 758.4500 371.7500 ;
        RECT 748.3000 369.7500 750.3000 371.7500 ;
        RECT 740.1500 369.7500 742.1500 371.7500 ;
        RECT 756.4500 376.8450 758.4500 378.8450 ;
        RECT 764.6000 376.8450 766.6000 378.8450 ;
        RECT 732.0000 398.1300 734.0000 400.1300 ;
        RECT 723.8500 398.1300 725.8500 400.1300 ;
        RECT 715.7000 398.1300 717.7000 400.1300 ;
        RECT 707.5500 398.1300 709.5500 400.1300 ;
        RECT 732.0000 391.0350 734.0000 393.0350 ;
        RECT 723.8500 391.0350 725.8500 393.0350 ;
        RECT 715.7000 391.0350 717.7000 393.0350 ;
        RECT 707.5500 391.0350 709.5500 393.0350 ;
        RECT 715.7000 412.3200 717.7000 414.3200 ;
        RECT 707.5500 412.3200 709.5500 414.3200 ;
        RECT 732.0000 405.2250 734.0000 407.2250 ;
        RECT 723.8500 405.2250 725.8500 407.2250 ;
        RECT 715.7000 405.2250 717.7000 407.2250 ;
        RECT 707.5500 405.2250 709.5500 407.2250 ;
        RECT 723.8500 412.3200 725.8500 414.3200 ;
        RECT 732.0000 412.3200 734.0000 414.3200 ;
        RECT 764.6000 398.1300 766.6000 400.1300 ;
        RECT 756.4500 398.1300 758.4500 400.1300 ;
        RECT 748.3000 398.1300 750.3000 400.1300 ;
        RECT 740.1500 398.1300 742.1500 400.1300 ;
        RECT 764.6000 391.0350 766.6000 393.0350 ;
        RECT 756.4500 391.0350 758.4500 393.0350 ;
        RECT 748.3000 391.0350 750.3000 393.0350 ;
        RECT 740.1500 391.0350 742.1500 393.0350 ;
        RECT 748.3000 412.3200 750.3000 414.3200 ;
        RECT 740.1500 412.3200 742.1500 414.3200 ;
        RECT 764.6000 405.2250 766.6000 407.2250 ;
        RECT 756.4500 405.2250 758.4500 407.2250 ;
        RECT 748.3000 405.2250 750.3000 407.2250 ;
        RECT 740.1500 405.2250 742.1500 407.2250 ;
        RECT 756.4500 412.3200 758.4500 414.3200 ;
        RECT 764.6000 412.3200 766.6000 414.3200 ;
        RECT 772.7500 383.9400 774.7500 385.9400 ;
        RECT 780.9000 383.9400 782.9000 385.9400 ;
        RECT 789.0500 383.9400 791.0500 385.9400 ;
        RECT 797.2000 383.9400 799.2000 385.9400 ;
        RECT 805.3500 383.9400 807.3500 385.9400 ;
        RECT 813.5000 383.9400 815.5000 385.9400 ;
        RECT 821.6500 383.9400 823.6500 385.9400 ;
        RECT 829.8000 383.9400 831.8000 385.9400 ;
        RECT 837.9500 383.9400 839.9500 385.9400 ;
        RECT 797.2000 362.6550 799.2000 364.6550 ;
        RECT 789.0500 362.6550 791.0500 364.6550 ;
        RECT 780.9000 362.6550 782.9000 364.6550 ;
        RECT 772.7500 362.6550 774.7500 364.6550 ;
        RECT 797.2000 355.5600 799.2000 357.5600 ;
        RECT 789.0500 355.5600 791.0500 357.5600 ;
        RECT 780.9000 355.5600 782.9000 357.5600 ;
        RECT 772.7500 355.5600 774.7500 357.5600 ;
        RECT 780.9000 376.8450 782.9000 378.8450 ;
        RECT 772.7500 376.8450 774.7500 378.8450 ;
        RECT 797.2000 369.7500 799.2000 371.7500 ;
        RECT 789.0500 369.7500 791.0500 371.7500 ;
        RECT 780.9000 369.7500 782.9000 371.7500 ;
        RECT 772.7500 369.7500 774.7500 371.7500 ;
        RECT 789.0500 376.8450 791.0500 378.8450 ;
        RECT 797.2000 376.8450 799.2000 378.8450 ;
        RECT 837.9500 362.6550 839.9500 364.6550 ;
        RECT 829.8000 362.6550 831.8000 364.6550 ;
        RECT 821.6500 362.6550 823.6500 364.6550 ;
        RECT 813.5000 362.6550 815.5000 364.6550 ;
        RECT 805.3500 362.6550 807.3500 364.6550 ;
        RECT 837.9500 355.5600 839.9500 357.5600 ;
        RECT 829.8000 355.5600 831.8000 357.5600 ;
        RECT 821.6500 355.5600 823.6500 357.5600 ;
        RECT 813.5000 355.5600 815.5000 357.5600 ;
        RECT 805.3500 355.5600 807.3500 357.5600 ;
        RECT 805.3500 369.7500 807.3500 371.7500 ;
        RECT 813.5000 369.7500 815.5000 371.7500 ;
        RECT 821.6500 369.7500 823.6500 371.7500 ;
        RECT 829.8000 369.7500 831.8000 371.7500 ;
        RECT 837.9500 369.7500 839.9500 371.7500 ;
        RECT 805.3500 376.8450 807.3500 378.8450 ;
        RECT 813.5000 376.8450 815.5000 378.8450 ;
        RECT 821.6500 376.8450 823.6500 378.8450 ;
        RECT 829.8000 376.8450 831.8000 378.8450 ;
        RECT 837.9500 376.8450 839.9500 378.8450 ;
        RECT 797.2000 398.1300 799.2000 400.1300 ;
        RECT 789.0500 398.1300 791.0500 400.1300 ;
        RECT 780.9000 398.1300 782.9000 400.1300 ;
        RECT 772.7500 398.1300 774.7500 400.1300 ;
        RECT 797.2000 391.0350 799.2000 393.0350 ;
        RECT 789.0500 391.0350 791.0500 393.0350 ;
        RECT 780.9000 391.0350 782.9000 393.0350 ;
        RECT 772.7500 391.0350 774.7500 393.0350 ;
        RECT 780.9000 412.3200 782.9000 414.3200 ;
        RECT 772.7500 412.3200 774.7500 414.3200 ;
        RECT 797.2000 405.2250 799.2000 407.2250 ;
        RECT 789.0500 405.2250 791.0500 407.2250 ;
        RECT 780.9000 405.2250 782.9000 407.2250 ;
        RECT 772.7500 405.2250 774.7500 407.2250 ;
        RECT 789.0500 412.3200 791.0500 414.3200 ;
        RECT 797.2000 412.3200 799.2000 414.3200 ;
        RECT 837.9500 398.1300 839.9500 400.1300 ;
        RECT 829.8000 398.1300 831.8000 400.1300 ;
        RECT 821.6500 398.1300 823.6500 400.1300 ;
        RECT 813.5000 398.1300 815.5000 400.1300 ;
        RECT 805.3500 398.1300 807.3500 400.1300 ;
        RECT 837.9500 391.0350 839.9500 393.0350 ;
        RECT 829.8000 391.0350 831.8000 393.0350 ;
        RECT 821.6500 391.0350 823.6500 393.0350 ;
        RECT 813.5000 391.0350 815.5000 393.0350 ;
        RECT 805.3500 391.0350 807.3500 393.0350 ;
        RECT 805.3500 405.2250 807.3500 407.2250 ;
        RECT 813.5000 405.2250 815.5000 407.2250 ;
        RECT 821.6500 405.2250 823.6500 407.2250 ;
        RECT 829.8000 405.2250 831.8000 407.2250 ;
        RECT 837.9500 405.2250 839.9500 407.2250 ;
        RECT 805.3500 412.3200 807.3500 414.3200 ;
        RECT 813.5000 412.3200 815.5000 414.3200 ;
        RECT 821.6500 412.3200 823.6500 414.3200 ;
        RECT 829.8000 412.3200 831.8000 414.3200 ;
        RECT 837.9500 412.3200 839.9500 414.3200 ;
        RECT 699.4000 483.2700 701.4000 485.2700 ;
        RECT 699.4000 476.1750 701.4000 478.1750 ;
        RECT 699.4000 469.0800 701.4000 471.0800 ;
        RECT 699.4000 461.9850 701.4000 463.9850 ;
        RECT 699.4000 454.8900 701.4000 456.8900 ;
        RECT 699.4000 447.7950 701.4000 449.7950 ;
        RECT 699.4000 440.7000 701.4000 442.7000 ;
        RECT 699.4000 433.6050 701.4000 435.6050 ;
        RECT 699.4000 426.5100 701.4000 428.5100 ;
        RECT 699.4000 497.4600 701.4000 499.4600 ;
        RECT 699.4000 490.3650 701.4000 492.3650 ;
        RECT 699.4000 504.5550 701.4000 506.5550 ;
        RECT 699.4000 511.6500 701.4000 513.6500 ;
        RECT 699.4000 518.7450 701.4000 520.7450 ;
        RECT 699.4000 525.8400 701.4000 527.8400 ;
        RECT 699.4000 532.9350 701.4000 534.9350 ;
        RECT 699.4000 540.0300 701.4000 542.0300 ;
        RECT 699.4000 547.1250 701.4000 549.1250 ;
        RECT 699.4000 554.2200 701.4000 556.2200 ;
        RECT 560.8500 454.8900 562.8500 456.8900 ;
        RECT 569.0000 454.8900 571.0000 456.8900 ;
        RECT 577.1500 454.8900 579.1500 456.8900 ;
        RECT 585.3000 454.8900 587.3000 456.8900 ;
        RECT 593.4500 454.8900 595.4500 456.8900 ;
        RECT 601.6000 454.8900 603.6000 456.8900 ;
        RECT 609.7500 454.8900 611.7500 456.8900 ;
        RECT 617.9000 454.8900 619.9000 456.8900 ;
        RECT 626.0500 454.8900 628.0500 456.8900 ;
        RECT 593.4500 426.5100 595.4500 428.5100 ;
        RECT 593.4500 433.6050 595.4500 435.6050 ;
        RECT 593.4500 440.7000 595.4500 442.7000 ;
        RECT 593.4500 447.7950 595.4500 449.7950 ;
        RECT 585.3000 433.6050 587.3000 435.6050 ;
        RECT 577.1500 433.6050 579.1500 435.6050 ;
        RECT 569.0000 433.6050 571.0000 435.6050 ;
        RECT 560.8500 433.6050 562.8500 435.6050 ;
        RECT 585.3000 426.5100 587.3000 428.5100 ;
        RECT 577.1500 426.5100 579.1500 428.5100 ;
        RECT 569.0000 426.5100 571.0000 428.5100 ;
        RECT 560.8500 426.5100 562.8500 428.5100 ;
        RECT 569.0000 447.7950 571.0000 449.7950 ;
        RECT 560.8500 447.7950 562.8500 449.7950 ;
        RECT 585.3000 440.7000 587.3000 442.7000 ;
        RECT 577.1500 440.7000 579.1500 442.7000 ;
        RECT 569.0000 440.7000 571.0000 442.7000 ;
        RECT 560.8500 440.7000 562.8500 442.7000 ;
        RECT 577.1500 447.7950 579.1500 449.7950 ;
        RECT 585.3000 447.7950 587.3000 449.7950 ;
        RECT 626.0500 433.6050 628.0500 435.6050 ;
        RECT 617.9000 433.6050 619.9000 435.6050 ;
        RECT 609.7500 433.6050 611.7500 435.6050 ;
        RECT 601.6000 433.6050 603.6000 435.6050 ;
        RECT 626.0500 426.5100 628.0500 428.5100 ;
        RECT 617.9000 426.5100 619.9000 428.5100 ;
        RECT 609.7500 426.5100 611.7500 428.5100 ;
        RECT 601.6000 426.5100 603.6000 428.5100 ;
        RECT 609.7500 447.7950 611.7500 449.7950 ;
        RECT 601.6000 447.7950 603.6000 449.7950 ;
        RECT 626.0500 440.7000 628.0500 442.7000 ;
        RECT 617.9000 440.7000 619.9000 442.7000 ;
        RECT 609.7500 440.7000 611.7500 442.7000 ;
        RECT 601.6000 440.7000 603.6000 442.7000 ;
        RECT 617.9000 447.7950 619.9000 449.7950 ;
        RECT 626.0500 447.7950 628.0500 449.7950 ;
        RECT 593.4500 461.9850 595.4500 463.9850 ;
        RECT 593.4500 469.0800 595.4500 471.0800 ;
        RECT 593.4500 476.1750 595.4500 478.1750 ;
        RECT 593.4500 483.2700 595.4500 485.2700 ;
        RECT 585.3000 469.0800 587.3000 471.0800 ;
        RECT 577.1500 469.0800 579.1500 471.0800 ;
        RECT 569.0000 469.0800 571.0000 471.0800 ;
        RECT 560.8500 469.0800 562.8500 471.0800 ;
        RECT 585.3000 461.9850 587.3000 463.9850 ;
        RECT 577.1500 461.9850 579.1500 463.9850 ;
        RECT 569.0000 461.9850 571.0000 463.9850 ;
        RECT 560.8500 461.9850 562.8500 463.9850 ;
        RECT 569.0000 483.2700 571.0000 485.2700 ;
        RECT 560.8500 483.2700 562.8500 485.2700 ;
        RECT 585.3000 476.1750 587.3000 478.1750 ;
        RECT 577.1500 476.1750 579.1500 478.1750 ;
        RECT 569.0000 476.1750 571.0000 478.1750 ;
        RECT 560.8500 476.1750 562.8500 478.1750 ;
        RECT 577.1500 483.2700 579.1500 485.2700 ;
        RECT 585.3000 483.2700 587.3000 485.2700 ;
        RECT 626.0500 469.0800 628.0500 471.0800 ;
        RECT 617.9000 469.0800 619.9000 471.0800 ;
        RECT 609.7500 469.0800 611.7500 471.0800 ;
        RECT 601.6000 469.0800 603.6000 471.0800 ;
        RECT 626.0500 461.9850 628.0500 463.9850 ;
        RECT 617.9000 461.9850 619.9000 463.9850 ;
        RECT 609.7500 461.9850 611.7500 463.9850 ;
        RECT 601.6000 461.9850 603.6000 463.9850 ;
        RECT 609.7500 483.2700 611.7500 485.2700 ;
        RECT 601.6000 483.2700 603.6000 485.2700 ;
        RECT 626.0500 476.1750 628.0500 478.1750 ;
        RECT 617.9000 476.1750 619.9000 478.1750 ;
        RECT 609.7500 476.1750 611.7500 478.1750 ;
        RECT 601.6000 476.1750 603.6000 478.1750 ;
        RECT 617.9000 483.2700 619.9000 485.2700 ;
        RECT 626.0500 483.2700 628.0500 485.2700 ;
        RECT 634.2000 454.8900 636.2000 456.8900 ;
        RECT 642.3500 454.8900 644.3500 456.8900 ;
        RECT 650.5000 454.8900 652.5000 456.8900 ;
        RECT 658.6500 454.8900 660.6500 456.8900 ;
        RECT 666.8000 454.8900 668.8000 456.8900 ;
        RECT 674.9500 454.8900 676.9500 456.8900 ;
        RECT 683.1000 454.8900 685.1000 456.8900 ;
        RECT 691.2500 454.8900 693.2500 456.8900 ;
        RECT 658.6500 433.6050 660.6500 435.6050 ;
        RECT 650.5000 433.6050 652.5000 435.6050 ;
        RECT 642.3500 433.6050 644.3500 435.6050 ;
        RECT 634.2000 433.6050 636.2000 435.6050 ;
        RECT 658.6500 426.5100 660.6500 428.5100 ;
        RECT 650.5000 426.5100 652.5000 428.5100 ;
        RECT 642.3500 426.5100 644.3500 428.5100 ;
        RECT 634.2000 426.5100 636.2000 428.5100 ;
        RECT 642.3500 447.7950 644.3500 449.7950 ;
        RECT 634.2000 447.7950 636.2000 449.7950 ;
        RECT 658.6500 440.7000 660.6500 442.7000 ;
        RECT 650.5000 440.7000 652.5000 442.7000 ;
        RECT 642.3500 440.7000 644.3500 442.7000 ;
        RECT 634.2000 440.7000 636.2000 442.7000 ;
        RECT 650.5000 447.7950 652.5000 449.7950 ;
        RECT 658.6500 447.7950 660.6500 449.7950 ;
        RECT 691.2500 433.6050 693.2500 435.6050 ;
        RECT 683.1000 433.6050 685.1000 435.6050 ;
        RECT 674.9500 433.6050 676.9500 435.6050 ;
        RECT 666.8000 433.6050 668.8000 435.6050 ;
        RECT 691.2500 426.5100 693.2500 428.5100 ;
        RECT 683.1000 426.5100 685.1000 428.5100 ;
        RECT 674.9500 426.5100 676.9500 428.5100 ;
        RECT 666.8000 426.5100 668.8000 428.5100 ;
        RECT 674.9500 447.7950 676.9500 449.7950 ;
        RECT 666.8000 447.7950 668.8000 449.7950 ;
        RECT 691.2500 440.7000 693.2500 442.7000 ;
        RECT 683.1000 440.7000 685.1000 442.7000 ;
        RECT 674.9500 440.7000 676.9500 442.7000 ;
        RECT 666.8000 440.7000 668.8000 442.7000 ;
        RECT 683.1000 447.7950 685.1000 449.7950 ;
        RECT 691.2500 447.7950 693.2500 449.7950 ;
        RECT 658.6500 469.0800 660.6500 471.0800 ;
        RECT 650.5000 469.0800 652.5000 471.0800 ;
        RECT 642.3500 469.0800 644.3500 471.0800 ;
        RECT 634.2000 469.0800 636.2000 471.0800 ;
        RECT 658.6500 461.9850 660.6500 463.9850 ;
        RECT 650.5000 461.9850 652.5000 463.9850 ;
        RECT 642.3500 461.9850 644.3500 463.9850 ;
        RECT 634.2000 461.9850 636.2000 463.9850 ;
        RECT 642.3500 483.2700 644.3500 485.2700 ;
        RECT 634.2000 483.2700 636.2000 485.2700 ;
        RECT 658.6500 476.1750 660.6500 478.1750 ;
        RECT 650.5000 476.1750 652.5000 478.1750 ;
        RECT 642.3500 476.1750 644.3500 478.1750 ;
        RECT 634.2000 476.1750 636.2000 478.1750 ;
        RECT 650.5000 483.2700 652.5000 485.2700 ;
        RECT 658.6500 483.2700 660.6500 485.2700 ;
        RECT 691.2500 469.0800 693.2500 471.0800 ;
        RECT 683.1000 469.0800 685.1000 471.0800 ;
        RECT 674.9500 469.0800 676.9500 471.0800 ;
        RECT 666.8000 469.0800 668.8000 471.0800 ;
        RECT 691.2500 461.9850 693.2500 463.9850 ;
        RECT 683.1000 461.9850 685.1000 463.9850 ;
        RECT 674.9500 461.9850 676.9500 463.9850 ;
        RECT 666.8000 461.9850 668.8000 463.9850 ;
        RECT 674.9500 483.2700 676.9500 485.2700 ;
        RECT 666.8000 483.2700 668.8000 485.2700 ;
        RECT 691.2500 476.1750 693.2500 478.1750 ;
        RECT 683.1000 476.1750 685.1000 478.1750 ;
        RECT 674.9500 476.1750 676.9500 478.1750 ;
        RECT 666.8000 476.1750 668.8000 478.1750 ;
        RECT 683.1000 483.2700 685.1000 485.2700 ;
        RECT 691.2500 483.2700 693.2500 485.2700 ;
        RECT 593.4500 490.3650 595.4500 492.3650 ;
        RECT 593.4500 497.4600 595.4500 499.4600 ;
        RECT 593.4500 504.5550 595.4500 506.5550 ;
        RECT 593.4500 511.6500 595.4500 513.6500 ;
        RECT 593.4500 518.7450 595.4500 520.7450 ;
        RECT 569.0000 504.5550 571.0000 506.5550 ;
        RECT 560.8500 504.5550 562.8500 506.5550 ;
        RECT 585.3000 497.4600 587.3000 499.4600 ;
        RECT 577.1500 497.4600 579.1500 499.4600 ;
        RECT 569.0000 497.4600 571.0000 499.4600 ;
        RECT 560.8500 497.4600 562.8500 499.4600 ;
        RECT 585.3000 490.3650 587.3000 492.3650 ;
        RECT 577.1500 490.3650 579.1500 492.3650 ;
        RECT 569.0000 490.3650 571.0000 492.3650 ;
        RECT 560.8500 490.3650 562.8500 492.3650 ;
        RECT 577.1500 504.5550 579.1500 506.5550 ;
        RECT 585.3000 504.5550 587.3000 506.5550 ;
        RECT 560.8500 511.6500 562.8500 513.6500 ;
        RECT 569.0000 511.6500 571.0000 513.6500 ;
        RECT 577.1500 511.6500 579.1500 513.6500 ;
        RECT 585.3000 511.6500 587.3000 513.6500 ;
        RECT 560.8500 518.7450 562.8500 520.7450 ;
        RECT 569.0000 518.7450 571.0000 520.7450 ;
        RECT 577.1500 518.7450 579.1500 520.7450 ;
        RECT 585.3000 518.7450 587.3000 520.7450 ;
        RECT 609.7500 504.5550 611.7500 506.5550 ;
        RECT 601.6000 504.5550 603.6000 506.5550 ;
        RECT 626.0500 497.4600 628.0500 499.4600 ;
        RECT 617.9000 497.4600 619.9000 499.4600 ;
        RECT 609.7500 497.4600 611.7500 499.4600 ;
        RECT 601.6000 497.4600 603.6000 499.4600 ;
        RECT 626.0500 490.3650 628.0500 492.3650 ;
        RECT 617.9000 490.3650 619.9000 492.3650 ;
        RECT 609.7500 490.3650 611.7500 492.3650 ;
        RECT 601.6000 490.3650 603.6000 492.3650 ;
        RECT 617.9000 504.5550 619.9000 506.5550 ;
        RECT 626.0500 504.5550 628.0500 506.5550 ;
        RECT 601.6000 511.6500 603.6000 513.6500 ;
        RECT 609.7500 511.6500 611.7500 513.6500 ;
        RECT 617.9000 511.6500 619.9000 513.6500 ;
        RECT 626.0500 511.6500 628.0500 513.6500 ;
        RECT 601.6000 518.7450 603.6000 520.7450 ;
        RECT 609.7500 518.7450 611.7500 520.7450 ;
        RECT 617.9000 518.7450 619.9000 520.7450 ;
        RECT 626.0500 518.7450 628.0500 520.7450 ;
        RECT 593.4500 525.8400 595.4500 527.8400 ;
        RECT 593.4500 532.9350 595.4500 534.9350 ;
        RECT 593.4500 540.0300 595.4500 542.0300 ;
        RECT 593.4500 547.1250 595.4500 549.1250 ;
        RECT 593.4500 554.2200 595.4500 556.2200 ;
        RECT 569.0000 540.0300 571.0000 542.0300 ;
        RECT 560.8500 540.0300 562.8500 542.0300 ;
        RECT 585.3000 532.9350 587.3000 534.9350 ;
        RECT 577.1500 532.9350 579.1500 534.9350 ;
        RECT 569.0000 532.9350 571.0000 534.9350 ;
        RECT 560.8500 532.9350 562.8500 534.9350 ;
        RECT 585.3000 525.8400 587.3000 527.8400 ;
        RECT 577.1500 525.8400 579.1500 527.8400 ;
        RECT 569.0000 525.8400 571.0000 527.8400 ;
        RECT 560.8500 525.8400 562.8500 527.8400 ;
        RECT 577.1500 540.0300 579.1500 542.0300 ;
        RECT 585.3000 540.0300 587.3000 542.0300 ;
        RECT 560.8500 547.1250 562.8500 549.1250 ;
        RECT 569.0000 547.1250 571.0000 549.1250 ;
        RECT 577.1500 547.1250 579.1500 549.1250 ;
        RECT 585.3000 547.1250 587.3000 549.1250 ;
        RECT 560.8500 554.2200 562.8500 556.2200 ;
        RECT 569.0000 554.2200 571.0000 556.2200 ;
        RECT 577.1500 554.2200 579.1500 556.2200 ;
        RECT 585.3000 554.2200 587.3000 556.2200 ;
        RECT 609.7500 540.0300 611.7500 542.0300 ;
        RECT 601.6000 540.0300 603.6000 542.0300 ;
        RECT 626.0500 532.9350 628.0500 534.9350 ;
        RECT 617.9000 532.9350 619.9000 534.9350 ;
        RECT 609.7500 532.9350 611.7500 534.9350 ;
        RECT 601.6000 532.9350 603.6000 534.9350 ;
        RECT 626.0500 525.8400 628.0500 527.8400 ;
        RECT 617.9000 525.8400 619.9000 527.8400 ;
        RECT 609.7500 525.8400 611.7500 527.8400 ;
        RECT 601.6000 525.8400 603.6000 527.8400 ;
        RECT 617.9000 540.0300 619.9000 542.0300 ;
        RECT 626.0500 540.0300 628.0500 542.0300 ;
        RECT 601.6000 547.1250 603.6000 549.1250 ;
        RECT 609.7500 547.1250 611.7500 549.1250 ;
        RECT 617.9000 547.1250 619.9000 549.1250 ;
        RECT 626.0500 547.1250 628.0500 549.1250 ;
        RECT 601.6000 554.2200 603.6000 556.2200 ;
        RECT 609.7500 554.2200 611.7500 556.2200 ;
        RECT 617.9000 554.2200 619.9000 556.2200 ;
        RECT 626.0500 554.2200 628.0500 556.2200 ;
        RECT 642.3500 504.5550 644.3500 506.5550 ;
        RECT 634.2000 504.5550 636.2000 506.5550 ;
        RECT 658.6500 497.4600 660.6500 499.4600 ;
        RECT 650.5000 497.4600 652.5000 499.4600 ;
        RECT 642.3500 497.4600 644.3500 499.4600 ;
        RECT 634.2000 497.4600 636.2000 499.4600 ;
        RECT 658.6500 490.3650 660.6500 492.3650 ;
        RECT 650.5000 490.3650 652.5000 492.3650 ;
        RECT 642.3500 490.3650 644.3500 492.3650 ;
        RECT 634.2000 490.3650 636.2000 492.3650 ;
        RECT 650.5000 504.5550 652.5000 506.5550 ;
        RECT 658.6500 504.5550 660.6500 506.5550 ;
        RECT 634.2000 511.6500 636.2000 513.6500 ;
        RECT 642.3500 511.6500 644.3500 513.6500 ;
        RECT 650.5000 511.6500 652.5000 513.6500 ;
        RECT 658.6500 511.6500 660.6500 513.6500 ;
        RECT 634.2000 518.7450 636.2000 520.7450 ;
        RECT 642.3500 518.7450 644.3500 520.7450 ;
        RECT 650.5000 518.7450 652.5000 520.7450 ;
        RECT 658.6500 518.7450 660.6500 520.7450 ;
        RECT 674.9500 504.5550 676.9500 506.5550 ;
        RECT 666.8000 504.5550 668.8000 506.5550 ;
        RECT 691.2500 497.4600 693.2500 499.4600 ;
        RECT 683.1000 497.4600 685.1000 499.4600 ;
        RECT 674.9500 497.4600 676.9500 499.4600 ;
        RECT 666.8000 497.4600 668.8000 499.4600 ;
        RECT 691.2500 490.3650 693.2500 492.3650 ;
        RECT 683.1000 490.3650 685.1000 492.3650 ;
        RECT 674.9500 490.3650 676.9500 492.3650 ;
        RECT 666.8000 490.3650 668.8000 492.3650 ;
        RECT 683.1000 504.5550 685.1000 506.5550 ;
        RECT 691.2500 504.5550 693.2500 506.5550 ;
        RECT 666.8000 511.6500 668.8000 513.6500 ;
        RECT 674.9500 511.6500 676.9500 513.6500 ;
        RECT 683.1000 511.6500 685.1000 513.6500 ;
        RECT 691.2500 511.6500 693.2500 513.6500 ;
        RECT 666.8000 518.7450 668.8000 520.7450 ;
        RECT 674.9500 518.7450 676.9500 520.7450 ;
        RECT 683.1000 518.7450 685.1000 520.7450 ;
        RECT 691.2500 518.7450 693.2500 520.7450 ;
        RECT 642.3500 540.0300 644.3500 542.0300 ;
        RECT 634.2000 540.0300 636.2000 542.0300 ;
        RECT 658.6500 532.9350 660.6500 534.9350 ;
        RECT 650.5000 532.9350 652.5000 534.9350 ;
        RECT 642.3500 532.9350 644.3500 534.9350 ;
        RECT 634.2000 532.9350 636.2000 534.9350 ;
        RECT 658.6500 525.8400 660.6500 527.8400 ;
        RECT 650.5000 525.8400 652.5000 527.8400 ;
        RECT 642.3500 525.8400 644.3500 527.8400 ;
        RECT 634.2000 525.8400 636.2000 527.8400 ;
        RECT 650.5000 540.0300 652.5000 542.0300 ;
        RECT 658.6500 540.0300 660.6500 542.0300 ;
        RECT 634.2000 547.1250 636.2000 549.1250 ;
        RECT 642.3500 547.1250 644.3500 549.1250 ;
        RECT 650.5000 547.1250 652.5000 549.1250 ;
        RECT 658.6500 547.1250 660.6500 549.1250 ;
        RECT 634.2000 554.2200 636.2000 556.2200 ;
        RECT 642.3500 554.2200 644.3500 556.2200 ;
        RECT 650.5000 554.2200 652.5000 556.2200 ;
        RECT 658.6500 554.2200 660.6500 556.2200 ;
        RECT 674.9500 540.0300 676.9500 542.0300 ;
        RECT 666.8000 540.0300 668.8000 542.0300 ;
        RECT 691.2500 532.9350 693.2500 534.9350 ;
        RECT 683.1000 532.9350 685.1000 534.9350 ;
        RECT 674.9500 532.9350 676.9500 534.9350 ;
        RECT 666.8000 532.9350 668.8000 534.9350 ;
        RECT 691.2500 525.8400 693.2500 527.8400 ;
        RECT 683.1000 525.8400 685.1000 527.8400 ;
        RECT 674.9500 525.8400 676.9500 527.8400 ;
        RECT 666.8000 525.8400 668.8000 527.8400 ;
        RECT 683.1000 540.0300 685.1000 542.0300 ;
        RECT 691.2500 540.0300 693.2500 542.0300 ;
        RECT 666.8000 547.1250 668.8000 549.1250 ;
        RECT 674.9500 547.1250 676.9500 549.1250 ;
        RECT 683.1000 547.1250 685.1000 549.1250 ;
        RECT 691.2500 547.1250 693.2500 549.1250 ;
        RECT 666.8000 554.2200 668.8000 556.2200 ;
        RECT 674.9500 554.2200 676.9500 556.2200 ;
        RECT 683.1000 554.2200 685.1000 556.2200 ;
        RECT 691.2500 554.2200 693.2500 556.2200 ;
        RECT 707.5500 454.8900 709.5500 456.8900 ;
        RECT 715.7000 454.8900 717.7000 456.8900 ;
        RECT 723.8500 454.8900 725.8500 456.8900 ;
        RECT 732.0000 454.8900 734.0000 456.8900 ;
        RECT 740.1500 454.8900 742.1500 456.8900 ;
        RECT 748.3000 454.8900 750.3000 456.8900 ;
        RECT 756.4500 454.8900 758.4500 456.8900 ;
        RECT 764.6000 454.8900 766.6000 456.8900 ;
        RECT 732.0000 433.6050 734.0000 435.6050 ;
        RECT 723.8500 433.6050 725.8500 435.6050 ;
        RECT 715.7000 433.6050 717.7000 435.6050 ;
        RECT 707.5500 433.6050 709.5500 435.6050 ;
        RECT 732.0000 426.5100 734.0000 428.5100 ;
        RECT 723.8500 426.5100 725.8500 428.5100 ;
        RECT 715.7000 426.5100 717.7000 428.5100 ;
        RECT 707.5500 426.5100 709.5500 428.5100 ;
        RECT 715.7000 447.7950 717.7000 449.7950 ;
        RECT 707.5500 447.7950 709.5500 449.7950 ;
        RECT 732.0000 440.7000 734.0000 442.7000 ;
        RECT 723.8500 440.7000 725.8500 442.7000 ;
        RECT 715.7000 440.7000 717.7000 442.7000 ;
        RECT 707.5500 440.7000 709.5500 442.7000 ;
        RECT 723.8500 447.7950 725.8500 449.7950 ;
        RECT 732.0000 447.7950 734.0000 449.7950 ;
        RECT 764.6000 433.6050 766.6000 435.6050 ;
        RECT 756.4500 433.6050 758.4500 435.6050 ;
        RECT 748.3000 433.6050 750.3000 435.6050 ;
        RECT 740.1500 433.6050 742.1500 435.6050 ;
        RECT 764.6000 426.5100 766.6000 428.5100 ;
        RECT 756.4500 426.5100 758.4500 428.5100 ;
        RECT 748.3000 426.5100 750.3000 428.5100 ;
        RECT 740.1500 426.5100 742.1500 428.5100 ;
        RECT 748.3000 447.7950 750.3000 449.7950 ;
        RECT 740.1500 447.7950 742.1500 449.7950 ;
        RECT 764.6000 440.7000 766.6000 442.7000 ;
        RECT 756.4500 440.7000 758.4500 442.7000 ;
        RECT 748.3000 440.7000 750.3000 442.7000 ;
        RECT 740.1500 440.7000 742.1500 442.7000 ;
        RECT 756.4500 447.7950 758.4500 449.7950 ;
        RECT 764.6000 447.7950 766.6000 449.7950 ;
        RECT 732.0000 469.0800 734.0000 471.0800 ;
        RECT 723.8500 469.0800 725.8500 471.0800 ;
        RECT 715.7000 469.0800 717.7000 471.0800 ;
        RECT 707.5500 469.0800 709.5500 471.0800 ;
        RECT 732.0000 461.9850 734.0000 463.9850 ;
        RECT 723.8500 461.9850 725.8500 463.9850 ;
        RECT 715.7000 461.9850 717.7000 463.9850 ;
        RECT 707.5500 461.9850 709.5500 463.9850 ;
        RECT 715.7000 483.2700 717.7000 485.2700 ;
        RECT 707.5500 483.2700 709.5500 485.2700 ;
        RECT 732.0000 476.1750 734.0000 478.1750 ;
        RECT 723.8500 476.1750 725.8500 478.1750 ;
        RECT 715.7000 476.1750 717.7000 478.1750 ;
        RECT 707.5500 476.1750 709.5500 478.1750 ;
        RECT 723.8500 483.2700 725.8500 485.2700 ;
        RECT 732.0000 483.2700 734.0000 485.2700 ;
        RECT 764.6000 469.0800 766.6000 471.0800 ;
        RECT 756.4500 469.0800 758.4500 471.0800 ;
        RECT 748.3000 469.0800 750.3000 471.0800 ;
        RECT 740.1500 469.0800 742.1500 471.0800 ;
        RECT 764.6000 461.9850 766.6000 463.9850 ;
        RECT 756.4500 461.9850 758.4500 463.9850 ;
        RECT 748.3000 461.9850 750.3000 463.9850 ;
        RECT 740.1500 461.9850 742.1500 463.9850 ;
        RECT 748.3000 483.2700 750.3000 485.2700 ;
        RECT 740.1500 483.2700 742.1500 485.2700 ;
        RECT 764.6000 476.1750 766.6000 478.1750 ;
        RECT 756.4500 476.1750 758.4500 478.1750 ;
        RECT 748.3000 476.1750 750.3000 478.1750 ;
        RECT 740.1500 476.1750 742.1500 478.1750 ;
        RECT 756.4500 483.2700 758.4500 485.2700 ;
        RECT 764.6000 483.2700 766.6000 485.2700 ;
        RECT 772.7500 454.8900 774.7500 456.8900 ;
        RECT 780.9000 454.8900 782.9000 456.8900 ;
        RECT 789.0500 454.8900 791.0500 456.8900 ;
        RECT 797.2000 454.8900 799.2000 456.8900 ;
        RECT 805.3500 454.8900 807.3500 456.8900 ;
        RECT 813.5000 454.8900 815.5000 456.8900 ;
        RECT 821.6500 454.8900 823.6500 456.8900 ;
        RECT 829.8000 454.8900 831.8000 456.8900 ;
        RECT 837.9500 454.8900 839.9500 456.8900 ;
        RECT 797.2000 433.6050 799.2000 435.6050 ;
        RECT 789.0500 433.6050 791.0500 435.6050 ;
        RECT 780.9000 433.6050 782.9000 435.6050 ;
        RECT 772.7500 433.6050 774.7500 435.6050 ;
        RECT 797.2000 426.5100 799.2000 428.5100 ;
        RECT 789.0500 426.5100 791.0500 428.5100 ;
        RECT 780.9000 426.5100 782.9000 428.5100 ;
        RECT 772.7500 426.5100 774.7500 428.5100 ;
        RECT 780.9000 447.7950 782.9000 449.7950 ;
        RECT 772.7500 447.7950 774.7500 449.7950 ;
        RECT 797.2000 440.7000 799.2000 442.7000 ;
        RECT 789.0500 440.7000 791.0500 442.7000 ;
        RECT 780.9000 440.7000 782.9000 442.7000 ;
        RECT 772.7500 440.7000 774.7500 442.7000 ;
        RECT 789.0500 447.7950 791.0500 449.7950 ;
        RECT 797.2000 447.7950 799.2000 449.7950 ;
        RECT 837.9500 433.6050 839.9500 435.6050 ;
        RECT 829.8000 433.6050 831.8000 435.6050 ;
        RECT 821.6500 433.6050 823.6500 435.6050 ;
        RECT 813.5000 433.6050 815.5000 435.6050 ;
        RECT 805.3500 433.6050 807.3500 435.6050 ;
        RECT 837.9500 426.5100 839.9500 428.5100 ;
        RECT 829.8000 426.5100 831.8000 428.5100 ;
        RECT 821.6500 426.5100 823.6500 428.5100 ;
        RECT 813.5000 426.5100 815.5000 428.5100 ;
        RECT 805.3500 426.5100 807.3500 428.5100 ;
        RECT 805.3500 440.7000 807.3500 442.7000 ;
        RECT 813.5000 440.7000 815.5000 442.7000 ;
        RECT 821.6500 440.7000 823.6500 442.7000 ;
        RECT 829.8000 440.7000 831.8000 442.7000 ;
        RECT 837.9500 440.7000 839.9500 442.7000 ;
        RECT 805.3500 447.7950 807.3500 449.7950 ;
        RECT 813.5000 447.7950 815.5000 449.7950 ;
        RECT 821.6500 447.7950 823.6500 449.7950 ;
        RECT 829.8000 447.7950 831.8000 449.7950 ;
        RECT 837.9500 447.7950 839.9500 449.7950 ;
        RECT 797.2000 469.0800 799.2000 471.0800 ;
        RECT 789.0500 469.0800 791.0500 471.0800 ;
        RECT 780.9000 469.0800 782.9000 471.0800 ;
        RECT 772.7500 469.0800 774.7500 471.0800 ;
        RECT 797.2000 461.9850 799.2000 463.9850 ;
        RECT 789.0500 461.9850 791.0500 463.9850 ;
        RECT 780.9000 461.9850 782.9000 463.9850 ;
        RECT 772.7500 461.9850 774.7500 463.9850 ;
        RECT 780.9000 483.2700 782.9000 485.2700 ;
        RECT 772.7500 483.2700 774.7500 485.2700 ;
        RECT 797.2000 476.1750 799.2000 478.1750 ;
        RECT 789.0500 476.1750 791.0500 478.1750 ;
        RECT 780.9000 476.1750 782.9000 478.1750 ;
        RECT 772.7500 476.1750 774.7500 478.1750 ;
        RECT 789.0500 483.2700 791.0500 485.2700 ;
        RECT 797.2000 483.2700 799.2000 485.2700 ;
        RECT 837.9500 469.0800 839.9500 471.0800 ;
        RECT 829.8000 469.0800 831.8000 471.0800 ;
        RECT 821.6500 469.0800 823.6500 471.0800 ;
        RECT 813.5000 469.0800 815.5000 471.0800 ;
        RECT 805.3500 469.0800 807.3500 471.0800 ;
        RECT 837.9500 461.9850 839.9500 463.9850 ;
        RECT 829.8000 461.9850 831.8000 463.9850 ;
        RECT 821.6500 461.9850 823.6500 463.9850 ;
        RECT 813.5000 461.9850 815.5000 463.9850 ;
        RECT 805.3500 461.9850 807.3500 463.9850 ;
        RECT 805.3500 476.1750 807.3500 478.1750 ;
        RECT 813.5000 476.1750 815.5000 478.1750 ;
        RECT 821.6500 476.1750 823.6500 478.1750 ;
        RECT 829.8000 476.1750 831.8000 478.1750 ;
        RECT 837.9500 476.1750 839.9500 478.1750 ;
        RECT 805.3500 483.2700 807.3500 485.2700 ;
        RECT 813.5000 483.2700 815.5000 485.2700 ;
        RECT 821.6500 483.2700 823.6500 485.2700 ;
        RECT 829.8000 483.2700 831.8000 485.2700 ;
        RECT 837.9500 483.2700 839.9500 485.2700 ;
        RECT 715.7000 504.5550 717.7000 506.5550 ;
        RECT 707.5500 504.5550 709.5500 506.5550 ;
        RECT 732.0000 497.4600 734.0000 499.4600 ;
        RECT 723.8500 497.4600 725.8500 499.4600 ;
        RECT 715.7000 497.4600 717.7000 499.4600 ;
        RECT 707.5500 497.4600 709.5500 499.4600 ;
        RECT 732.0000 490.3650 734.0000 492.3650 ;
        RECT 723.8500 490.3650 725.8500 492.3650 ;
        RECT 715.7000 490.3650 717.7000 492.3650 ;
        RECT 707.5500 490.3650 709.5500 492.3650 ;
        RECT 723.8500 504.5550 725.8500 506.5550 ;
        RECT 732.0000 504.5550 734.0000 506.5550 ;
        RECT 707.5500 511.6500 709.5500 513.6500 ;
        RECT 715.7000 511.6500 717.7000 513.6500 ;
        RECT 723.8500 511.6500 725.8500 513.6500 ;
        RECT 732.0000 511.6500 734.0000 513.6500 ;
        RECT 707.5500 518.7450 709.5500 520.7450 ;
        RECT 715.7000 518.7450 717.7000 520.7450 ;
        RECT 723.8500 518.7450 725.8500 520.7450 ;
        RECT 732.0000 518.7450 734.0000 520.7450 ;
        RECT 748.3000 504.5550 750.3000 506.5550 ;
        RECT 740.1500 504.5550 742.1500 506.5550 ;
        RECT 764.6000 497.4600 766.6000 499.4600 ;
        RECT 756.4500 497.4600 758.4500 499.4600 ;
        RECT 748.3000 497.4600 750.3000 499.4600 ;
        RECT 740.1500 497.4600 742.1500 499.4600 ;
        RECT 764.6000 490.3650 766.6000 492.3650 ;
        RECT 756.4500 490.3650 758.4500 492.3650 ;
        RECT 748.3000 490.3650 750.3000 492.3650 ;
        RECT 740.1500 490.3650 742.1500 492.3650 ;
        RECT 756.4500 504.5550 758.4500 506.5550 ;
        RECT 764.6000 504.5550 766.6000 506.5550 ;
        RECT 740.1500 511.6500 742.1500 513.6500 ;
        RECT 748.3000 511.6500 750.3000 513.6500 ;
        RECT 756.4500 511.6500 758.4500 513.6500 ;
        RECT 764.6000 511.6500 766.6000 513.6500 ;
        RECT 740.1500 518.7450 742.1500 520.7450 ;
        RECT 748.3000 518.7450 750.3000 520.7450 ;
        RECT 756.4500 518.7450 758.4500 520.7450 ;
        RECT 764.6000 518.7450 766.6000 520.7450 ;
        RECT 715.7000 540.0300 717.7000 542.0300 ;
        RECT 707.5500 540.0300 709.5500 542.0300 ;
        RECT 732.0000 532.9350 734.0000 534.9350 ;
        RECT 723.8500 532.9350 725.8500 534.9350 ;
        RECT 715.7000 532.9350 717.7000 534.9350 ;
        RECT 707.5500 532.9350 709.5500 534.9350 ;
        RECT 732.0000 525.8400 734.0000 527.8400 ;
        RECT 723.8500 525.8400 725.8500 527.8400 ;
        RECT 715.7000 525.8400 717.7000 527.8400 ;
        RECT 707.5500 525.8400 709.5500 527.8400 ;
        RECT 723.8500 540.0300 725.8500 542.0300 ;
        RECT 732.0000 540.0300 734.0000 542.0300 ;
        RECT 707.5500 547.1250 709.5500 549.1250 ;
        RECT 715.7000 547.1250 717.7000 549.1250 ;
        RECT 723.8500 547.1250 725.8500 549.1250 ;
        RECT 732.0000 547.1250 734.0000 549.1250 ;
        RECT 707.5500 554.2200 709.5500 556.2200 ;
        RECT 715.7000 554.2200 717.7000 556.2200 ;
        RECT 723.8500 554.2200 725.8500 556.2200 ;
        RECT 732.0000 554.2200 734.0000 556.2200 ;
        RECT 748.3000 540.0300 750.3000 542.0300 ;
        RECT 740.1500 540.0300 742.1500 542.0300 ;
        RECT 764.6000 532.9350 766.6000 534.9350 ;
        RECT 756.4500 532.9350 758.4500 534.9350 ;
        RECT 748.3000 532.9350 750.3000 534.9350 ;
        RECT 740.1500 532.9350 742.1500 534.9350 ;
        RECT 764.6000 525.8400 766.6000 527.8400 ;
        RECT 756.4500 525.8400 758.4500 527.8400 ;
        RECT 748.3000 525.8400 750.3000 527.8400 ;
        RECT 740.1500 525.8400 742.1500 527.8400 ;
        RECT 756.4500 540.0300 758.4500 542.0300 ;
        RECT 764.6000 540.0300 766.6000 542.0300 ;
        RECT 740.1500 547.1250 742.1500 549.1250 ;
        RECT 748.3000 547.1250 750.3000 549.1250 ;
        RECT 756.4500 547.1250 758.4500 549.1250 ;
        RECT 764.6000 547.1250 766.6000 549.1250 ;
        RECT 740.1500 554.2200 742.1500 556.2200 ;
        RECT 748.3000 554.2200 750.3000 556.2200 ;
        RECT 756.4500 554.2200 758.4500 556.2200 ;
        RECT 764.6000 554.2200 766.6000 556.2200 ;
        RECT 780.9000 504.5550 782.9000 506.5550 ;
        RECT 772.7500 504.5550 774.7500 506.5550 ;
        RECT 797.2000 497.4600 799.2000 499.4600 ;
        RECT 789.0500 497.4600 791.0500 499.4600 ;
        RECT 780.9000 497.4600 782.9000 499.4600 ;
        RECT 772.7500 497.4600 774.7500 499.4600 ;
        RECT 797.2000 490.3650 799.2000 492.3650 ;
        RECT 789.0500 490.3650 791.0500 492.3650 ;
        RECT 780.9000 490.3650 782.9000 492.3650 ;
        RECT 772.7500 490.3650 774.7500 492.3650 ;
        RECT 789.0500 504.5550 791.0500 506.5550 ;
        RECT 797.2000 504.5550 799.2000 506.5550 ;
        RECT 772.7500 511.6500 774.7500 513.6500 ;
        RECT 780.9000 511.6500 782.9000 513.6500 ;
        RECT 789.0500 511.6500 791.0500 513.6500 ;
        RECT 797.2000 511.6500 799.2000 513.6500 ;
        RECT 772.7500 518.7450 774.7500 520.7450 ;
        RECT 780.9000 518.7450 782.9000 520.7450 ;
        RECT 789.0500 518.7450 791.0500 520.7450 ;
        RECT 797.2000 518.7450 799.2000 520.7450 ;
        RECT 821.6500 490.3650 823.6500 492.3650 ;
        RECT 821.6500 497.4600 823.6500 499.4600 ;
        RECT 821.6500 504.5550 823.6500 506.5550 ;
        RECT 813.5000 504.5550 815.5000 506.5550 ;
        RECT 805.3500 504.5550 807.3500 506.5550 ;
        RECT 813.5000 497.4600 815.5000 499.4600 ;
        RECT 805.3500 497.4600 807.3500 499.4600 ;
        RECT 805.3500 490.3650 807.3500 492.3650 ;
        RECT 813.5000 490.3650 815.5000 492.3650 ;
        RECT 837.9500 504.5550 839.9500 506.5550 ;
        RECT 829.8000 504.5550 831.8000 506.5550 ;
        RECT 837.9500 497.4600 839.9500 499.4600 ;
        RECT 829.8000 497.4600 831.8000 499.4600 ;
        RECT 829.8000 490.3650 831.8000 492.3650 ;
        RECT 837.9500 490.3650 839.9500 492.3650 ;
        RECT 805.3500 511.6500 807.3500 513.6500 ;
        RECT 813.5000 511.6500 815.5000 513.6500 ;
        RECT 821.6500 511.6500 823.6500 513.6500 ;
        RECT 829.8000 511.6500 831.8000 513.6500 ;
        RECT 837.9500 511.6500 839.9500 513.6500 ;
        RECT 805.3500 518.7450 807.3500 520.7450 ;
        RECT 813.5000 518.7450 815.5000 520.7450 ;
        RECT 821.6500 518.7450 823.6500 520.7450 ;
        RECT 829.8000 518.7450 831.8000 520.7450 ;
        RECT 837.9500 518.7450 839.9500 520.7450 ;
        RECT 780.9000 540.0300 782.9000 542.0300 ;
        RECT 772.7500 540.0300 774.7500 542.0300 ;
        RECT 797.2000 532.9350 799.2000 534.9350 ;
        RECT 789.0500 532.9350 791.0500 534.9350 ;
        RECT 780.9000 532.9350 782.9000 534.9350 ;
        RECT 772.7500 532.9350 774.7500 534.9350 ;
        RECT 797.2000 525.8400 799.2000 527.8400 ;
        RECT 789.0500 525.8400 791.0500 527.8400 ;
        RECT 780.9000 525.8400 782.9000 527.8400 ;
        RECT 772.7500 525.8400 774.7500 527.8400 ;
        RECT 789.0500 540.0300 791.0500 542.0300 ;
        RECT 797.2000 540.0300 799.2000 542.0300 ;
        RECT 772.7500 547.1250 774.7500 549.1250 ;
        RECT 780.9000 547.1250 782.9000 549.1250 ;
        RECT 789.0500 547.1250 791.0500 549.1250 ;
        RECT 797.2000 547.1250 799.2000 549.1250 ;
        RECT 772.7500 554.2200 774.7500 556.2200 ;
        RECT 780.9000 554.2200 782.9000 556.2200 ;
        RECT 789.0500 554.2200 791.0500 556.2200 ;
        RECT 797.2000 554.2200 799.2000 556.2200 ;
        RECT 821.6500 525.8400 823.6500 527.8400 ;
        RECT 821.6500 532.9350 823.6500 534.9350 ;
        RECT 821.6500 540.0300 823.6500 542.0300 ;
        RECT 813.5000 540.0300 815.5000 542.0300 ;
        RECT 805.3500 540.0300 807.3500 542.0300 ;
        RECT 813.5000 532.9350 815.5000 534.9350 ;
        RECT 805.3500 532.9350 807.3500 534.9350 ;
        RECT 805.3500 525.8400 807.3500 527.8400 ;
        RECT 813.5000 525.8400 815.5000 527.8400 ;
        RECT 837.9500 540.0300 839.9500 542.0300 ;
        RECT 829.8000 540.0300 831.8000 542.0300 ;
        RECT 837.9500 532.9350 839.9500 534.9350 ;
        RECT 829.8000 532.9350 831.8000 534.9350 ;
        RECT 829.8000 525.8400 831.8000 527.8400 ;
        RECT 837.9500 525.8400 839.9500 527.8400 ;
        RECT 805.3500 547.1250 807.3500 549.1250 ;
        RECT 813.5000 547.1250 815.5000 549.1250 ;
        RECT 821.6500 547.1250 823.6500 549.1250 ;
        RECT 829.8000 547.1250 831.8000 549.1250 ;
        RECT 837.9500 547.1250 839.9500 549.1250 ;
        RECT 805.3500 554.2200 807.3500 556.2200 ;
        RECT 813.5000 554.2200 815.5000 556.2200 ;
        RECT 821.6500 554.2200 823.6500 556.2200 ;
        RECT 829.8000 554.2200 831.8000 556.2200 ;
        RECT 837.9500 554.2200 839.9500 556.2200 ;
        RECT 903.1500 419.4150 905.1500 421.4150 ;
        RECT 895.0000 419.4150 897.0000 421.4150 ;
        RECT 886.8500 419.4150 888.8500 421.4150 ;
        RECT 878.7000 419.4150 880.7000 421.4150 ;
        RECT 870.5500 419.4150 872.5500 421.4150 ;
        RECT 862.4000 419.4150 864.4000 421.4150 ;
        RECT 854.2500 419.4150 856.2500 421.4150 ;
        RECT 846.1000 419.4150 848.1000 421.4150 ;
        RECT 943.9000 419.4150 945.9000 421.4150 ;
        RECT 935.7500 419.4150 937.7500 421.4150 ;
        RECT 927.6000 419.4150 929.6000 421.4150 ;
        RECT 919.4500 419.4150 921.4500 421.4150 ;
        RECT 911.3000 419.4150 913.3000 421.4150 ;
        RECT 952.0500 419.4150 954.0500 421.4150 ;
        RECT 960.2000 419.4150 962.2000 421.4150 ;
        RECT 968.3500 419.4150 970.3500 421.4150 ;
        RECT 976.5000 419.4150 978.5000 421.4150 ;
        RECT 1112.0000 419.4150 1114.0000 421.4150 ;
        RECT 1074.0000 419.4150 1076.0000 421.4150 ;
        RECT 984.6500 419.4150 986.6500 421.4150 ;
        RECT 992.8000 419.4150 994.8000 421.4150 ;
        RECT 1000.9500 419.4150 1002.9500 421.4150 ;
        RECT 1009.1000 419.4150 1011.1000 421.4150 ;
        RECT 1017.2500 419.4150 1019.2500 421.4150 ;
        RECT 1025.4000 419.4150 1027.4000 421.4150 ;
        RECT 1033.5500 419.4150 1035.5500 421.4150 ;
        RECT 1041.7000 419.4150 1043.7000 421.4150 ;
        RECT 1049.8500 419.4150 1051.8500 421.4150 ;
        RECT 1058.0000 419.4150 1060.0000 421.4150 ;
        RECT 903.1500 348.4650 905.1500 350.4650 ;
        RECT 895.0000 348.4650 897.0000 350.4650 ;
        RECT 886.8500 348.4650 888.8500 350.4650 ;
        RECT 878.7000 348.4650 880.7000 350.4650 ;
        RECT 870.5500 348.4650 872.5500 350.4650 ;
        RECT 862.4000 348.4650 864.4000 350.4650 ;
        RECT 854.2500 348.4650 856.2500 350.4650 ;
        RECT 846.1000 348.4650 848.1000 350.4650 ;
        RECT 943.9000 348.4650 945.9000 350.4650 ;
        RECT 935.7500 348.4650 937.7500 350.4650 ;
        RECT 927.6000 348.4650 929.6000 350.4650 ;
        RECT 919.4500 348.4650 921.4500 350.4650 ;
        RECT 911.3000 348.4650 913.3000 350.4650 ;
        RECT 952.0500 348.4650 954.0500 350.4650 ;
        RECT 960.2000 348.4650 962.2000 350.4650 ;
        RECT 968.3500 348.4650 970.3500 350.4650 ;
        RECT 976.5000 348.4650 978.5000 350.4650 ;
        RECT 870.5500 291.7050 872.5500 293.7050 ;
        RECT 862.4000 291.7050 864.4000 293.7050 ;
        RECT 854.2500 291.7050 856.2500 293.7050 ;
        RECT 846.1000 291.7050 848.1000 293.7050 ;
        RECT 870.5500 284.6100 872.5500 286.6100 ;
        RECT 862.4000 284.6100 864.4000 286.6100 ;
        RECT 854.2500 284.6100 856.2500 286.6100 ;
        RECT 846.1000 284.6100 848.1000 286.6100 ;
        RECT 854.2500 298.8000 856.2500 300.8000 ;
        RECT 846.1000 298.8000 848.1000 300.8000 ;
        RECT 862.4000 298.8000 864.4000 300.8000 ;
        RECT 870.5500 298.8000 872.5500 300.8000 ;
        RECT 846.1000 305.8950 848.1000 307.8950 ;
        RECT 854.2500 305.8950 856.2500 307.8950 ;
        RECT 862.4000 305.8950 864.4000 307.8950 ;
        RECT 870.5500 305.8950 872.5500 307.8950 ;
        RECT 846.1000 312.9900 848.1000 314.9900 ;
        RECT 854.2500 312.9900 856.2500 314.9900 ;
        RECT 862.4000 312.9900 864.4000 314.9900 ;
        RECT 870.5500 312.9900 872.5500 314.9900 ;
        RECT 903.1500 291.7050 905.1500 293.7050 ;
        RECT 895.0000 291.7050 897.0000 293.7050 ;
        RECT 886.8500 291.7050 888.8500 293.7050 ;
        RECT 878.7000 291.7050 880.7000 293.7050 ;
        RECT 903.1500 284.6100 905.1500 286.6100 ;
        RECT 895.0000 284.6100 897.0000 286.6100 ;
        RECT 886.8500 284.6100 888.8500 286.6100 ;
        RECT 878.7000 284.6100 880.7000 286.6100 ;
        RECT 886.8500 298.8000 888.8500 300.8000 ;
        RECT 878.7000 298.8000 880.7000 300.8000 ;
        RECT 895.0000 298.8000 897.0000 300.8000 ;
        RECT 903.1500 298.8000 905.1500 300.8000 ;
        RECT 878.7000 305.8950 880.7000 307.8950 ;
        RECT 886.8500 305.8950 888.8500 307.8950 ;
        RECT 895.0000 305.8950 897.0000 307.8950 ;
        RECT 903.1500 305.8950 905.1500 307.8950 ;
        RECT 878.7000 312.9900 880.7000 314.9900 ;
        RECT 886.8500 312.9900 888.8500 314.9900 ;
        RECT 895.0000 312.9900 897.0000 314.9900 ;
        RECT 903.1500 312.9900 905.1500 314.9900 ;
        RECT 870.5500 327.1800 872.5500 329.1800 ;
        RECT 862.4000 327.1800 864.4000 329.1800 ;
        RECT 854.2500 327.1800 856.2500 329.1800 ;
        RECT 846.1000 327.1800 848.1000 329.1800 ;
        RECT 870.5500 320.0850 872.5500 322.0850 ;
        RECT 862.4000 320.0850 864.4000 322.0850 ;
        RECT 854.2500 320.0850 856.2500 322.0850 ;
        RECT 846.1000 320.0850 848.1000 322.0850 ;
        RECT 854.2500 341.3700 856.2500 343.3700 ;
        RECT 846.1000 341.3700 848.1000 343.3700 ;
        RECT 870.5500 334.2750 872.5500 336.2750 ;
        RECT 862.4000 334.2750 864.4000 336.2750 ;
        RECT 854.2500 334.2750 856.2500 336.2750 ;
        RECT 846.1000 334.2750 848.1000 336.2750 ;
        RECT 862.4000 341.3700 864.4000 343.3700 ;
        RECT 870.5500 341.3700 872.5500 343.3700 ;
        RECT 903.1500 327.1800 905.1500 329.1800 ;
        RECT 895.0000 327.1800 897.0000 329.1800 ;
        RECT 886.8500 327.1800 888.8500 329.1800 ;
        RECT 878.7000 327.1800 880.7000 329.1800 ;
        RECT 903.1500 320.0850 905.1500 322.0850 ;
        RECT 895.0000 320.0850 897.0000 322.0850 ;
        RECT 886.8500 320.0850 888.8500 322.0850 ;
        RECT 878.7000 320.0850 880.7000 322.0850 ;
        RECT 886.8500 341.3700 888.8500 343.3700 ;
        RECT 878.7000 341.3700 880.7000 343.3700 ;
        RECT 903.1500 334.2750 905.1500 336.2750 ;
        RECT 895.0000 334.2750 897.0000 336.2750 ;
        RECT 886.8500 334.2750 888.8500 336.2750 ;
        RECT 878.7000 334.2750 880.7000 336.2750 ;
        RECT 895.0000 341.3700 897.0000 343.3700 ;
        RECT 903.1500 341.3700 905.1500 343.3700 ;
        RECT 943.9000 284.6100 945.9000 286.6100 ;
        RECT 943.9000 291.7050 945.9000 293.7050 ;
        RECT 943.9000 298.8000 945.9000 300.8000 ;
        RECT 943.9000 305.8950 945.9000 307.8950 ;
        RECT 943.9000 312.9900 945.9000 314.9900 ;
        RECT 935.7500 291.7050 937.7500 293.7050 ;
        RECT 927.6000 291.7050 929.6000 293.7050 ;
        RECT 919.4500 291.7050 921.4500 293.7050 ;
        RECT 911.3000 291.7050 913.3000 293.7050 ;
        RECT 935.7500 284.6100 937.7500 286.6100 ;
        RECT 927.6000 284.6100 929.6000 286.6100 ;
        RECT 919.4500 284.6100 921.4500 286.6100 ;
        RECT 911.3000 284.6100 913.3000 286.6100 ;
        RECT 919.4500 298.8000 921.4500 300.8000 ;
        RECT 911.3000 298.8000 913.3000 300.8000 ;
        RECT 927.6000 298.8000 929.6000 300.8000 ;
        RECT 935.7500 298.8000 937.7500 300.8000 ;
        RECT 911.3000 305.8950 913.3000 307.8950 ;
        RECT 919.4500 305.8950 921.4500 307.8950 ;
        RECT 927.6000 305.8950 929.6000 307.8950 ;
        RECT 935.7500 305.8950 937.7500 307.8950 ;
        RECT 911.3000 312.9900 913.3000 314.9900 ;
        RECT 919.4500 312.9900 921.4500 314.9900 ;
        RECT 927.6000 312.9900 929.6000 314.9900 ;
        RECT 935.7500 312.9900 937.7500 314.9900 ;
        RECT 976.5000 291.7050 978.5000 293.7050 ;
        RECT 968.3500 291.7050 970.3500 293.7050 ;
        RECT 960.2000 291.7050 962.2000 293.7050 ;
        RECT 952.0500 291.7050 954.0500 293.7050 ;
        RECT 976.5000 284.6100 978.5000 286.6100 ;
        RECT 968.3500 284.6100 970.3500 286.6100 ;
        RECT 960.2000 284.6100 962.2000 286.6100 ;
        RECT 952.0500 284.6100 954.0500 286.6100 ;
        RECT 960.2000 298.8000 962.2000 300.8000 ;
        RECT 952.0500 298.8000 954.0500 300.8000 ;
        RECT 968.3500 298.8000 970.3500 300.8000 ;
        RECT 976.5000 298.8000 978.5000 300.8000 ;
        RECT 952.0500 305.8950 954.0500 307.8950 ;
        RECT 960.2000 305.8950 962.2000 307.8950 ;
        RECT 968.3500 305.8950 970.3500 307.8950 ;
        RECT 976.5000 305.8950 978.5000 307.8950 ;
        RECT 952.0500 312.9900 954.0500 314.9900 ;
        RECT 960.2000 312.9900 962.2000 314.9900 ;
        RECT 968.3500 312.9900 970.3500 314.9900 ;
        RECT 976.5000 312.9900 978.5000 314.9900 ;
        RECT 943.9000 320.0850 945.9000 322.0850 ;
        RECT 943.9000 327.1800 945.9000 329.1800 ;
        RECT 943.9000 334.2750 945.9000 336.2750 ;
        RECT 943.9000 341.3700 945.9000 343.3700 ;
        RECT 935.7500 327.1800 937.7500 329.1800 ;
        RECT 927.6000 327.1800 929.6000 329.1800 ;
        RECT 919.4500 327.1800 921.4500 329.1800 ;
        RECT 911.3000 327.1800 913.3000 329.1800 ;
        RECT 935.7500 320.0850 937.7500 322.0850 ;
        RECT 927.6000 320.0850 929.6000 322.0850 ;
        RECT 919.4500 320.0850 921.4500 322.0850 ;
        RECT 911.3000 320.0850 913.3000 322.0850 ;
        RECT 919.4500 341.3700 921.4500 343.3700 ;
        RECT 911.3000 341.3700 913.3000 343.3700 ;
        RECT 935.7500 334.2750 937.7500 336.2750 ;
        RECT 927.6000 334.2750 929.6000 336.2750 ;
        RECT 919.4500 334.2750 921.4500 336.2750 ;
        RECT 911.3000 334.2750 913.3000 336.2750 ;
        RECT 927.6000 341.3700 929.6000 343.3700 ;
        RECT 935.7500 341.3700 937.7500 343.3700 ;
        RECT 976.5000 327.1800 978.5000 329.1800 ;
        RECT 968.3500 327.1800 970.3500 329.1800 ;
        RECT 960.2000 327.1800 962.2000 329.1800 ;
        RECT 952.0500 327.1800 954.0500 329.1800 ;
        RECT 976.5000 320.0850 978.5000 322.0850 ;
        RECT 968.3500 320.0850 970.3500 322.0850 ;
        RECT 960.2000 320.0850 962.2000 322.0850 ;
        RECT 952.0500 320.0850 954.0500 322.0850 ;
        RECT 960.2000 341.3700 962.2000 343.3700 ;
        RECT 952.0500 341.3700 954.0500 343.3700 ;
        RECT 976.5000 334.2750 978.5000 336.2750 ;
        RECT 968.3500 334.2750 970.3500 336.2750 ;
        RECT 960.2000 334.2750 962.2000 336.2750 ;
        RECT 952.0500 334.2750 954.0500 336.2750 ;
        RECT 968.3500 341.3700 970.3500 343.3700 ;
        RECT 976.5000 341.3700 978.5000 343.3700 ;
        RECT 846.1000 383.9400 848.1000 385.9400 ;
        RECT 854.2500 383.9400 856.2500 385.9400 ;
        RECT 862.4000 383.9400 864.4000 385.9400 ;
        RECT 870.5500 383.9400 872.5500 385.9400 ;
        RECT 878.7000 383.9400 880.7000 385.9400 ;
        RECT 886.8500 383.9400 888.8500 385.9400 ;
        RECT 895.0000 383.9400 897.0000 385.9400 ;
        RECT 903.1500 383.9400 905.1500 385.9400 ;
        RECT 870.5500 362.6550 872.5500 364.6550 ;
        RECT 862.4000 362.6550 864.4000 364.6550 ;
        RECT 854.2500 362.6550 856.2500 364.6550 ;
        RECT 846.1000 362.6550 848.1000 364.6550 ;
        RECT 870.5500 355.5600 872.5500 357.5600 ;
        RECT 862.4000 355.5600 864.4000 357.5600 ;
        RECT 854.2500 355.5600 856.2500 357.5600 ;
        RECT 846.1000 355.5600 848.1000 357.5600 ;
        RECT 854.2500 376.8450 856.2500 378.8450 ;
        RECT 846.1000 376.8450 848.1000 378.8450 ;
        RECT 870.5500 369.7500 872.5500 371.7500 ;
        RECT 862.4000 369.7500 864.4000 371.7500 ;
        RECT 854.2500 369.7500 856.2500 371.7500 ;
        RECT 846.1000 369.7500 848.1000 371.7500 ;
        RECT 862.4000 376.8450 864.4000 378.8450 ;
        RECT 870.5500 376.8450 872.5500 378.8450 ;
        RECT 903.1500 362.6550 905.1500 364.6550 ;
        RECT 895.0000 362.6550 897.0000 364.6550 ;
        RECT 886.8500 362.6550 888.8500 364.6550 ;
        RECT 878.7000 362.6550 880.7000 364.6550 ;
        RECT 903.1500 355.5600 905.1500 357.5600 ;
        RECT 895.0000 355.5600 897.0000 357.5600 ;
        RECT 886.8500 355.5600 888.8500 357.5600 ;
        RECT 878.7000 355.5600 880.7000 357.5600 ;
        RECT 886.8500 376.8450 888.8500 378.8450 ;
        RECT 878.7000 376.8450 880.7000 378.8450 ;
        RECT 903.1500 369.7500 905.1500 371.7500 ;
        RECT 895.0000 369.7500 897.0000 371.7500 ;
        RECT 886.8500 369.7500 888.8500 371.7500 ;
        RECT 878.7000 369.7500 880.7000 371.7500 ;
        RECT 895.0000 376.8450 897.0000 378.8450 ;
        RECT 903.1500 376.8450 905.1500 378.8450 ;
        RECT 870.5500 398.1300 872.5500 400.1300 ;
        RECT 862.4000 398.1300 864.4000 400.1300 ;
        RECT 854.2500 398.1300 856.2500 400.1300 ;
        RECT 846.1000 398.1300 848.1000 400.1300 ;
        RECT 870.5500 391.0350 872.5500 393.0350 ;
        RECT 862.4000 391.0350 864.4000 393.0350 ;
        RECT 854.2500 391.0350 856.2500 393.0350 ;
        RECT 846.1000 391.0350 848.1000 393.0350 ;
        RECT 854.2500 412.3200 856.2500 414.3200 ;
        RECT 846.1000 412.3200 848.1000 414.3200 ;
        RECT 870.5500 405.2250 872.5500 407.2250 ;
        RECT 862.4000 405.2250 864.4000 407.2250 ;
        RECT 854.2500 405.2250 856.2500 407.2250 ;
        RECT 846.1000 405.2250 848.1000 407.2250 ;
        RECT 862.4000 412.3200 864.4000 414.3200 ;
        RECT 870.5500 412.3200 872.5500 414.3200 ;
        RECT 903.1500 398.1300 905.1500 400.1300 ;
        RECT 895.0000 398.1300 897.0000 400.1300 ;
        RECT 886.8500 398.1300 888.8500 400.1300 ;
        RECT 878.7000 398.1300 880.7000 400.1300 ;
        RECT 903.1500 391.0350 905.1500 393.0350 ;
        RECT 895.0000 391.0350 897.0000 393.0350 ;
        RECT 886.8500 391.0350 888.8500 393.0350 ;
        RECT 878.7000 391.0350 880.7000 393.0350 ;
        RECT 886.8500 412.3200 888.8500 414.3200 ;
        RECT 878.7000 412.3200 880.7000 414.3200 ;
        RECT 903.1500 405.2250 905.1500 407.2250 ;
        RECT 895.0000 405.2250 897.0000 407.2250 ;
        RECT 886.8500 405.2250 888.8500 407.2250 ;
        RECT 878.7000 405.2250 880.7000 407.2250 ;
        RECT 895.0000 412.3200 897.0000 414.3200 ;
        RECT 903.1500 412.3200 905.1500 414.3200 ;
        RECT 911.3000 383.9400 913.3000 385.9400 ;
        RECT 919.4500 383.9400 921.4500 385.9400 ;
        RECT 927.6000 383.9400 929.6000 385.9400 ;
        RECT 935.7500 383.9400 937.7500 385.9400 ;
        RECT 943.9000 383.9400 945.9000 385.9400 ;
        RECT 952.0500 383.9400 954.0500 385.9400 ;
        RECT 960.2000 383.9400 962.2000 385.9400 ;
        RECT 968.3500 383.9400 970.3500 385.9400 ;
        RECT 976.5000 383.9400 978.5000 385.9400 ;
        RECT 943.9000 355.5600 945.9000 357.5600 ;
        RECT 943.9000 362.6550 945.9000 364.6550 ;
        RECT 943.9000 369.7500 945.9000 371.7500 ;
        RECT 943.9000 376.8450 945.9000 378.8450 ;
        RECT 935.7500 362.6550 937.7500 364.6550 ;
        RECT 927.6000 362.6550 929.6000 364.6550 ;
        RECT 919.4500 362.6550 921.4500 364.6550 ;
        RECT 911.3000 362.6550 913.3000 364.6550 ;
        RECT 935.7500 355.5600 937.7500 357.5600 ;
        RECT 927.6000 355.5600 929.6000 357.5600 ;
        RECT 919.4500 355.5600 921.4500 357.5600 ;
        RECT 911.3000 355.5600 913.3000 357.5600 ;
        RECT 919.4500 376.8450 921.4500 378.8450 ;
        RECT 911.3000 376.8450 913.3000 378.8450 ;
        RECT 935.7500 369.7500 937.7500 371.7500 ;
        RECT 927.6000 369.7500 929.6000 371.7500 ;
        RECT 919.4500 369.7500 921.4500 371.7500 ;
        RECT 911.3000 369.7500 913.3000 371.7500 ;
        RECT 927.6000 376.8450 929.6000 378.8450 ;
        RECT 935.7500 376.8450 937.7500 378.8450 ;
        RECT 976.5000 362.6550 978.5000 364.6550 ;
        RECT 968.3500 362.6550 970.3500 364.6550 ;
        RECT 960.2000 362.6550 962.2000 364.6550 ;
        RECT 952.0500 362.6550 954.0500 364.6550 ;
        RECT 976.5000 355.5600 978.5000 357.5600 ;
        RECT 968.3500 355.5600 970.3500 357.5600 ;
        RECT 960.2000 355.5600 962.2000 357.5600 ;
        RECT 952.0500 355.5600 954.0500 357.5600 ;
        RECT 960.2000 376.8450 962.2000 378.8450 ;
        RECT 952.0500 376.8450 954.0500 378.8450 ;
        RECT 976.5000 369.7500 978.5000 371.7500 ;
        RECT 968.3500 369.7500 970.3500 371.7500 ;
        RECT 960.2000 369.7500 962.2000 371.7500 ;
        RECT 952.0500 369.7500 954.0500 371.7500 ;
        RECT 968.3500 376.8450 970.3500 378.8450 ;
        RECT 976.5000 376.8450 978.5000 378.8450 ;
        RECT 943.9000 391.0350 945.9000 393.0350 ;
        RECT 943.9000 398.1300 945.9000 400.1300 ;
        RECT 943.9000 405.2250 945.9000 407.2250 ;
        RECT 943.9000 412.3200 945.9000 414.3200 ;
        RECT 935.7500 398.1300 937.7500 400.1300 ;
        RECT 927.6000 398.1300 929.6000 400.1300 ;
        RECT 919.4500 398.1300 921.4500 400.1300 ;
        RECT 911.3000 398.1300 913.3000 400.1300 ;
        RECT 935.7500 391.0350 937.7500 393.0350 ;
        RECT 927.6000 391.0350 929.6000 393.0350 ;
        RECT 919.4500 391.0350 921.4500 393.0350 ;
        RECT 911.3000 391.0350 913.3000 393.0350 ;
        RECT 919.4500 412.3200 921.4500 414.3200 ;
        RECT 911.3000 412.3200 913.3000 414.3200 ;
        RECT 935.7500 405.2250 937.7500 407.2250 ;
        RECT 927.6000 405.2250 929.6000 407.2250 ;
        RECT 919.4500 405.2250 921.4500 407.2250 ;
        RECT 911.3000 405.2250 913.3000 407.2250 ;
        RECT 927.6000 412.3200 929.6000 414.3200 ;
        RECT 935.7500 412.3200 937.7500 414.3200 ;
        RECT 976.5000 398.1300 978.5000 400.1300 ;
        RECT 968.3500 398.1300 970.3500 400.1300 ;
        RECT 960.2000 398.1300 962.2000 400.1300 ;
        RECT 952.0500 398.1300 954.0500 400.1300 ;
        RECT 976.5000 391.0350 978.5000 393.0350 ;
        RECT 968.3500 391.0350 970.3500 393.0350 ;
        RECT 960.2000 391.0350 962.2000 393.0350 ;
        RECT 952.0500 391.0350 954.0500 393.0350 ;
        RECT 960.2000 412.3200 962.2000 414.3200 ;
        RECT 952.0500 412.3200 954.0500 414.3200 ;
        RECT 976.5000 405.2250 978.5000 407.2250 ;
        RECT 968.3500 405.2250 970.3500 407.2250 ;
        RECT 960.2000 405.2250 962.2000 407.2250 ;
        RECT 952.0500 405.2250 954.0500 407.2250 ;
        RECT 968.3500 412.3200 970.3500 414.3200 ;
        RECT 976.5000 412.3200 978.5000 414.3200 ;
        RECT 1074.0000 348.4650 1076.0000 350.4650 ;
        RECT 1112.0000 348.4650 1114.0000 350.4650 ;
        RECT 984.6500 348.4650 986.6500 350.4650 ;
        RECT 992.8000 348.4650 994.8000 350.4650 ;
        RECT 1000.9500 348.4650 1002.9500 350.4650 ;
        RECT 1009.1000 348.4650 1011.1000 350.4650 ;
        RECT 1017.2500 348.4650 1019.2500 350.4650 ;
        RECT 1025.4000 348.4650 1027.4000 350.4650 ;
        RECT 1033.5500 348.4650 1035.5500 350.4650 ;
        RECT 1041.7000 348.4650 1043.7000 350.4650 ;
        RECT 1049.8500 348.4650 1051.8500 350.4650 ;
        RECT 1058.0000 348.4650 1060.0000 350.4650 ;
        RECT 1049.8500 284.6100 1051.8500 286.6100 ;
        RECT 1049.8500 291.7050 1051.8500 293.7050 ;
        RECT 1049.8500 298.8000 1051.8500 300.8000 ;
        RECT 1049.8500 305.8950 1051.8500 307.8950 ;
        RECT 1049.8500 312.9900 1051.8500 314.9900 ;
        RECT 1049.8500 320.0850 1051.8500 322.0850 ;
        RECT 1049.8500 327.1800 1051.8500 329.1800 ;
        RECT 1049.8500 334.2750 1051.8500 336.2750 ;
        RECT 1049.8500 341.3700 1051.8500 343.3700 ;
        RECT 1009.1000 291.7050 1011.1000 293.7050 ;
        RECT 1000.9500 291.7050 1002.9500 293.7050 ;
        RECT 992.8000 291.7050 994.8000 293.7050 ;
        RECT 984.6500 291.7050 986.6500 293.7050 ;
        RECT 1009.1000 284.6100 1011.1000 286.6100 ;
        RECT 1000.9500 284.6100 1002.9500 286.6100 ;
        RECT 992.8000 284.6100 994.8000 286.6100 ;
        RECT 984.6500 284.6100 986.6500 286.6100 ;
        RECT 992.8000 298.8000 994.8000 300.8000 ;
        RECT 984.6500 298.8000 986.6500 300.8000 ;
        RECT 1000.9500 298.8000 1002.9500 300.8000 ;
        RECT 1009.1000 298.8000 1011.1000 300.8000 ;
        RECT 984.6500 305.8950 986.6500 307.8950 ;
        RECT 992.8000 305.8950 994.8000 307.8950 ;
        RECT 1000.9500 305.8950 1002.9500 307.8950 ;
        RECT 1009.1000 305.8950 1011.1000 307.8950 ;
        RECT 984.6500 312.9900 986.6500 314.9900 ;
        RECT 992.8000 312.9900 994.8000 314.9900 ;
        RECT 1000.9500 312.9900 1002.9500 314.9900 ;
        RECT 1009.1000 312.9900 1011.1000 314.9900 ;
        RECT 1041.7000 291.7050 1043.7000 293.7050 ;
        RECT 1033.5500 291.7050 1035.5500 293.7050 ;
        RECT 1025.4000 291.7050 1027.4000 293.7050 ;
        RECT 1017.2500 291.7050 1019.2500 293.7050 ;
        RECT 1041.7000 284.6100 1043.7000 286.6100 ;
        RECT 1033.5500 284.6100 1035.5500 286.6100 ;
        RECT 1025.4000 284.6100 1027.4000 286.6100 ;
        RECT 1017.2500 284.6100 1019.2500 286.6100 ;
        RECT 1025.4000 298.8000 1027.4000 300.8000 ;
        RECT 1017.2500 298.8000 1019.2500 300.8000 ;
        RECT 1033.5500 298.8000 1035.5500 300.8000 ;
        RECT 1041.7000 298.8000 1043.7000 300.8000 ;
        RECT 1017.2500 305.8950 1019.2500 307.8950 ;
        RECT 1025.4000 305.8950 1027.4000 307.8950 ;
        RECT 1033.5500 305.8950 1035.5500 307.8950 ;
        RECT 1041.7000 305.8950 1043.7000 307.8950 ;
        RECT 1017.2500 312.9900 1019.2500 314.9900 ;
        RECT 1025.4000 312.9900 1027.4000 314.9900 ;
        RECT 1033.5500 312.9900 1035.5500 314.9900 ;
        RECT 1041.7000 312.9900 1043.7000 314.9900 ;
        RECT 1009.1000 327.1800 1011.1000 329.1800 ;
        RECT 1000.9500 327.1800 1002.9500 329.1800 ;
        RECT 992.8000 327.1800 994.8000 329.1800 ;
        RECT 984.6500 327.1800 986.6500 329.1800 ;
        RECT 1009.1000 320.0850 1011.1000 322.0850 ;
        RECT 1000.9500 320.0850 1002.9500 322.0850 ;
        RECT 992.8000 320.0850 994.8000 322.0850 ;
        RECT 984.6500 320.0850 986.6500 322.0850 ;
        RECT 992.8000 341.3700 994.8000 343.3700 ;
        RECT 984.6500 341.3700 986.6500 343.3700 ;
        RECT 1009.1000 334.2750 1011.1000 336.2750 ;
        RECT 1000.9500 334.2750 1002.9500 336.2750 ;
        RECT 992.8000 334.2750 994.8000 336.2750 ;
        RECT 984.6500 334.2750 986.6500 336.2750 ;
        RECT 1000.9500 341.3700 1002.9500 343.3700 ;
        RECT 1009.1000 341.3700 1011.1000 343.3700 ;
        RECT 1041.7000 327.1800 1043.7000 329.1800 ;
        RECT 1033.5500 327.1800 1035.5500 329.1800 ;
        RECT 1025.4000 327.1800 1027.4000 329.1800 ;
        RECT 1017.2500 327.1800 1019.2500 329.1800 ;
        RECT 1041.7000 320.0850 1043.7000 322.0850 ;
        RECT 1033.5500 320.0850 1035.5500 322.0850 ;
        RECT 1025.4000 320.0850 1027.4000 322.0850 ;
        RECT 1017.2500 320.0850 1019.2500 322.0850 ;
        RECT 1025.4000 341.3700 1027.4000 343.3700 ;
        RECT 1017.2500 341.3700 1019.2500 343.3700 ;
        RECT 1041.7000 334.2750 1043.7000 336.2750 ;
        RECT 1033.5500 334.2750 1035.5500 336.2750 ;
        RECT 1025.4000 334.2750 1027.4000 336.2750 ;
        RECT 1017.2500 334.2750 1019.2500 336.2750 ;
        RECT 1033.5500 341.3700 1035.5500 343.3700 ;
        RECT 1041.7000 341.3700 1043.7000 343.3700 ;
        RECT 1058.0000 291.7050 1060.0000 293.7050 ;
        RECT 1058.0000 284.6100 1060.0000 286.6100 ;
        RECT 1074.0000 291.7050 1076.0000 293.7050 ;
        RECT 1074.0000 284.6100 1076.0000 286.6100 ;
        RECT 1058.0000 298.8000 1060.0000 300.8000 ;
        RECT 1058.0000 305.8950 1060.0000 307.8950 ;
        RECT 1058.0000 312.9900 1060.0000 314.9900 ;
        RECT 1074.0000 305.8950 1076.0000 307.8950 ;
        RECT 1074.0000 298.8000 1076.0000 300.8000 ;
        RECT 1074.0000 312.9900 1076.0000 314.9900 ;
        RECT 1112.0000 284.6100 1114.0000 286.6100 ;
        RECT 1112.0000 291.7050 1114.0000 293.7050 ;
        RECT 1112.0000 305.8950 1114.0000 307.8950 ;
        RECT 1112.0000 298.8000 1114.0000 300.8000 ;
        RECT 1112.0000 312.9900 1114.0000 314.9900 ;
        RECT 1058.0000 327.1800 1060.0000 329.1800 ;
        RECT 1058.0000 320.0850 1060.0000 322.0850 ;
        RECT 1074.0000 320.0850 1076.0000 322.0850 ;
        RECT 1074.0000 327.1800 1076.0000 329.1800 ;
        RECT 1058.0000 341.3700 1060.0000 343.3700 ;
        RECT 1058.0000 334.2750 1060.0000 336.2750 ;
        RECT 1074.0000 341.3700 1076.0000 343.3700 ;
        RECT 1074.0000 334.2750 1076.0000 336.2750 ;
        RECT 1112.0000 320.0850 1114.0000 322.0850 ;
        RECT 1112.0000 327.1800 1114.0000 329.1800 ;
        RECT 1112.0000 334.2750 1114.0000 336.2750 ;
        RECT 1112.0000 341.3700 1114.0000 343.3700 ;
        RECT 1049.8500 355.5600 1051.8500 357.5600 ;
        RECT 1049.8500 362.6550 1051.8500 364.6550 ;
        RECT 1049.8500 369.7500 1051.8500 371.7500 ;
        RECT 1049.8500 376.8450 1051.8500 378.8450 ;
        RECT 1049.8500 383.9400 1051.8500 385.9400 ;
        RECT 1049.8500 391.0350 1051.8500 393.0350 ;
        RECT 1049.8500 398.1300 1051.8500 400.1300 ;
        RECT 1049.8500 405.2250 1051.8500 407.2250 ;
        RECT 1049.8500 412.3200 1051.8500 414.3200 ;
        RECT 984.6500 383.9400 986.6500 385.9400 ;
        RECT 992.8000 383.9400 994.8000 385.9400 ;
        RECT 1000.9500 383.9400 1002.9500 385.9400 ;
        RECT 1009.1000 383.9400 1011.1000 385.9400 ;
        RECT 1017.2500 383.9400 1019.2500 385.9400 ;
        RECT 1025.4000 383.9400 1027.4000 385.9400 ;
        RECT 1033.5500 383.9400 1035.5500 385.9400 ;
        RECT 1041.7000 383.9400 1043.7000 385.9400 ;
        RECT 1009.1000 362.6550 1011.1000 364.6550 ;
        RECT 1000.9500 362.6550 1002.9500 364.6550 ;
        RECT 992.8000 362.6550 994.8000 364.6550 ;
        RECT 984.6500 362.6550 986.6500 364.6550 ;
        RECT 1009.1000 355.5600 1011.1000 357.5600 ;
        RECT 1000.9500 355.5600 1002.9500 357.5600 ;
        RECT 992.8000 355.5600 994.8000 357.5600 ;
        RECT 984.6500 355.5600 986.6500 357.5600 ;
        RECT 992.8000 376.8450 994.8000 378.8450 ;
        RECT 984.6500 376.8450 986.6500 378.8450 ;
        RECT 1009.1000 369.7500 1011.1000 371.7500 ;
        RECT 1000.9500 369.7500 1002.9500 371.7500 ;
        RECT 992.8000 369.7500 994.8000 371.7500 ;
        RECT 984.6500 369.7500 986.6500 371.7500 ;
        RECT 1000.9500 376.8450 1002.9500 378.8450 ;
        RECT 1009.1000 376.8450 1011.1000 378.8450 ;
        RECT 1041.7000 362.6550 1043.7000 364.6550 ;
        RECT 1033.5500 362.6550 1035.5500 364.6550 ;
        RECT 1025.4000 362.6550 1027.4000 364.6550 ;
        RECT 1017.2500 362.6550 1019.2500 364.6550 ;
        RECT 1041.7000 355.5600 1043.7000 357.5600 ;
        RECT 1033.5500 355.5600 1035.5500 357.5600 ;
        RECT 1025.4000 355.5600 1027.4000 357.5600 ;
        RECT 1017.2500 355.5600 1019.2500 357.5600 ;
        RECT 1025.4000 376.8450 1027.4000 378.8450 ;
        RECT 1017.2500 376.8450 1019.2500 378.8450 ;
        RECT 1041.7000 369.7500 1043.7000 371.7500 ;
        RECT 1033.5500 369.7500 1035.5500 371.7500 ;
        RECT 1025.4000 369.7500 1027.4000 371.7500 ;
        RECT 1017.2500 369.7500 1019.2500 371.7500 ;
        RECT 1033.5500 376.8450 1035.5500 378.8450 ;
        RECT 1041.7000 376.8450 1043.7000 378.8450 ;
        RECT 1009.1000 398.1300 1011.1000 400.1300 ;
        RECT 1000.9500 398.1300 1002.9500 400.1300 ;
        RECT 992.8000 398.1300 994.8000 400.1300 ;
        RECT 984.6500 398.1300 986.6500 400.1300 ;
        RECT 1009.1000 391.0350 1011.1000 393.0350 ;
        RECT 1000.9500 391.0350 1002.9500 393.0350 ;
        RECT 992.8000 391.0350 994.8000 393.0350 ;
        RECT 984.6500 391.0350 986.6500 393.0350 ;
        RECT 992.8000 412.3200 994.8000 414.3200 ;
        RECT 984.6500 412.3200 986.6500 414.3200 ;
        RECT 1009.1000 405.2250 1011.1000 407.2250 ;
        RECT 1000.9500 405.2250 1002.9500 407.2250 ;
        RECT 992.8000 405.2250 994.8000 407.2250 ;
        RECT 984.6500 405.2250 986.6500 407.2250 ;
        RECT 1000.9500 412.3200 1002.9500 414.3200 ;
        RECT 1009.1000 412.3200 1011.1000 414.3200 ;
        RECT 1041.7000 398.1300 1043.7000 400.1300 ;
        RECT 1033.5500 398.1300 1035.5500 400.1300 ;
        RECT 1025.4000 398.1300 1027.4000 400.1300 ;
        RECT 1017.2500 398.1300 1019.2500 400.1300 ;
        RECT 1041.7000 391.0350 1043.7000 393.0350 ;
        RECT 1033.5500 391.0350 1035.5500 393.0350 ;
        RECT 1025.4000 391.0350 1027.4000 393.0350 ;
        RECT 1017.2500 391.0350 1019.2500 393.0350 ;
        RECT 1025.4000 412.3200 1027.4000 414.3200 ;
        RECT 1017.2500 412.3200 1019.2500 414.3200 ;
        RECT 1041.7000 405.2250 1043.7000 407.2250 ;
        RECT 1033.5500 405.2250 1035.5500 407.2250 ;
        RECT 1025.4000 405.2250 1027.4000 407.2250 ;
        RECT 1017.2500 405.2250 1019.2500 407.2250 ;
        RECT 1033.5500 412.3200 1035.5500 414.3200 ;
        RECT 1041.7000 412.3200 1043.7000 414.3200 ;
        RECT 1074.0000 383.9400 1076.0000 385.9400 ;
        RECT 1112.0000 383.9400 1114.0000 385.9400 ;
        RECT 1058.0000 383.9400 1060.0000 385.9400 ;
        RECT 1058.0000 362.6550 1060.0000 364.6550 ;
        RECT 1058.0000 355.5600 1060.0000 357.5600 ;
        RECT 1074.0000 355.5600 1076.0000 357.5600 ;
        RECT 1074.0000 362.6550 1076.0000 364.6550 ;
        RECT 1058.0000 369.7500 1060.0000 371.7500 ;
        RECT 1058.0000 376.8450 1060.0000 378.8450 ;
        RECT 1074.0000 369.7500 1076.0000 371.7500 ;
        RECT 1074.0000 376.8450 1076.0000 378.8450 ;
        RECT 1112.0000 355.5600 1114.0000 357.5600 ;
        RECT 1112.0000 362.6550 1114.0000 364.6550 ;
        RECT 1112.0000 369.7500 1114.0000 371.7500 ;
        RECT 1112.0000 376.8450 1114.0000 378.8450 ;
        RECT 1058.0000 398.1300 1060.0000 400.1300 ;
        RECT 1058.0000 391.0350 1060.0000 393.0350 ;
        RECT 1074.0000 398.1300 1076.0000 400.1300 ;
        RECT 1074.0000 391.0350 1076.0000 393.0350 ;
        RECT 1058.0000 412.3200 1060.0000 414.3200 ;
        RECT 1058.0000 405.2250 1060.0000 407.2250 ;
        RECT 1074.0000 412.3200 1076.0000 414.3200 ;
        RECT 1074.0000 405.2250 1076.0000 407.2250 ;
        RECT 1112.0000 391.0350 1114.0000 393.0350 ;
        RECT 1112.0000 398.1300 1114.0000 400.1300 ;
        RECT 1112.0000 405.2250 1114.0000 407.2250 ;
        RECT 1112.0000 412.3200 1114.0000 414.3200 ;
        RECT 846.1000 454.8900 848.1000 456.8900 ;
        RECT 854.2500 454.8900 856.2500 456.8900 ;
        RECT 862.4000 454.8900 864.4000 456.8900 ;
        RECT 870.5500 454.8900 872.5500 456.8900 ;
        RECT 878.7000 454.8900 880.7000 456.8900 ;
        RECT 886.8500 454.8900 888.8500 456.8900 ;
        RECT 895.0000 454.8900 897.0000 456.8900 ;
        RECT 903.1500 454.8900 905.1500 456.8900 ;
        RECT 870.5500 433.6050 872.5500 435.6050 ;
        RECT 862.4000 433.6050 864.4000 435.6050 ;
        RECT 854.2500 433.6050 856.2500 435.6050 ;
        RECT 846.1000 433.6050 848.1000 435.6050 ;
        RECT 870.5500 426.5100 872.5500 428.5100 ;
        RECT 862.4000 426.5100 864.4000 428.5100 ;
        RECT 854.2500 426.5100 856.2500 428.5100 ;
        RECT 846.1000 426.5100 848.1000 428.5100 ;
        RECT 854.2500 447.7950 856.2500 449.7950 ;
        RECT 846.1000 447.7950 848.1000 449.7950 ;
        RECT 870.5500 440.7000 872.5500 442.7000 ;
        RECT 862.4000 440.7000 864.4000 442.7000 ;
        RECT 854.2500 440.7000 856.2500 442.7000 ;
        RECT 846.1000 440.7000 848.1000 442.7000 ;
        RECT 862.4000 447.7950 864.4000 449.7950 ;
        RECT 870.5500 447.7950 872.5500 449.7950 ;
        RECT 903.1500 433.6050 905.1500 435.6050 ;
        RECT 895.0000 433.6050 897.0000 435.6050 ;
        RECT 886.8500 433.6050 888.8500 435.6050 ;
        RECT 878.7000 433.6050 880.7000 435.6050 ;
        RECT 903.1500 426.5100 905.1500 428.5100 ;
        RECT 895.0000 426.5100 897.0000 428.5100 ;
        RECT 886.8500 426.5100 888.8500 428.5100 ;
        RECT 878.7000 426.5100 880.7000 428.5100 ;
        RECT 886.8500 447.7950 888.8500 449.7950 ;
        RECT 878.7000 447.7950 880.7000 449.7950 ;
        RECT 903.1500 440.7000 905.1500 442.7000 ;
        RECT 895.0000 440.7000 897.0000 442.7000 ;
        RECT 886.8500 440.7000 888.8500 442.7000 ;
        RECT 878.7000 440.7000 880.7000 442.7000 ;
        RECT 895.0000 447.7950 897.0000 449.7950 ;
        RECT 903.1500 447.7950 905.1500 449.7950 ;
        RECT 870.5500 469.0800 872.5500 471.0800 ;
        RECT 862.4000 469.0800 864.4000 471.0800 ;
        RECT 854.2500 469.0800 856.2500 471.0800 ;
        RECT 846.1000 469.0800 848.1000 471.0800 ;
        RECT 870.5500 461.9850 872.5500 463.9850 ;
        RECT 862.4000 461.9850 864.4000 463.9850 ;
        RECT 854.2500 461.9850 856.2500 463.9850 ;
        RECT 846.1000 461.9850 848.1000 463.9850 ;
        RECT 854.2500 483.2700 856.2500 485.2700 ;
        RECT 846.1000 483.2700 848.1000 485.2700 ;
        RECT 870.5500 476.1750 872.5500 478.1750 ;
        RECT 862.4000 476.1750 864.4000 478.1750 ;
        RECT 854.2500 476.1750 856.2500 478.1750 ;
        RECT 846.1000 476.1750 848.1000 478.1750 ;
        RECT 862.4000 483.2700 864.4000 485.2700 ;
        RECT 870.5500 483.2700 872.5500 485.2700 ;
        RECT 903.1500 469.0800 905.1500 471.0800 ;
        RECT 895.0000 469.0800 897.0000 471.0800 ;
        RECT 886.8500 469.0800 888.8500 471.0800 ;
        RECT 878.7000 469.0800 880.7000 471.0800 ;
        RECT 903.1500 461.9850 905.1500 463.9850 ;
        RECT 895.0000 461.9850 897.0000 463.9850 ;
        RECT 886.8500 461.9850 888.8500 463.9850 ;
        RECT 878.7000 461.9850 880.7000 463.9850 ;
        RECT 886.8500 483.2700 888.8500 485.2700 ;
        RECT 878.7000 483.2700 880.7000 485.2700 ;
        RECT 903.1500 476.1750 905.1500 478.1750 ;
        RECT 895.0000 476.1750 897.0000 478.1750 ;
        RECT 886.8500 476.1750 888.8500 478.1750 ;
        RECT 878.7000 476.1750 880.7000 478.1750 ;
        RECT 895.0000 483.2700 897.0000 485.2700 ;
        RECT 903.1500 483.2700 905.1500 485.2700 ;
        RECT 911.3000 454.8900 913.3000 456.8900 ;
        RECT 919.4500 454.8900 921.4500 456.8900 ;
        RECT 927.6000 454.8900 929.6000 456.8900 ;
        RECT 935.7500 454.8900 937.7500 456.8900 ;
        RECT 943.9000 454.8900 945.9000 456.8900 ;
        RECT 952.0500 454.8900 954.0500 456.8900 ;
        RECT 960.2000 454.8900 962.2000 456.8900 ;
        RECT 968.3500 454.8900 970.3500 456.8900 ;
        RECT 976.5000 454.8900 978.5000 456.8900 ;
        RECT 943.9000 426.5100 945.9000 428.5100 ;
        RECT 943.9000 433.6050 945.9000 435.6050 ;
        RECT 943.9000 440.7000 945.9000 442.7000 ;
        RECT 943.9000 447.7950 945.9000 449.7950 ;
        RECT 935.7500 433.6050 937.7500 435.6050 ;
        RECT 927.6000 433.6050 929.6000 435.6050 ;
        RECT 919.4500 433.6050 921.4500 435.6050 ;
        RECT 911.3000 433.6050 913.3000 435.6050 ;
        RECT 935.7500 426.5100 937.7500 428.5100 ;
        RECT 927.6000 426.5100 929.6000 428.5100 ;
        RECT 919.4500 426.5100 921.4500 428.5100 ;
        RECT 911.3000 426.5100 913.3000 428.5100 ;
        RECT 919.4500 447.7950 921.4500 449.7950 ;
        RECT 911.3000 447.7950 913.3000 449.7950 ;
        RECT 935.7500 440.7000 937.7500 442.7000 ;
        RECT 927.6000 440.7000 929.6000 442.7000 ;
        RECT 919.4500 440.7000 921.4500 442.7000 ;
        RECT 911.3000 440.7000 913.3000 442.7000 ;
        RECT 927.6000 447.7950 929.6000 449.7950 ;
        RECT 935.7500 447.7950 937.7500 449.7950 ;
        RECT 976.5000 433.6050 978.5000 435.6050 ;
        RECT 968.3500 433.6050 970.3500 435.6050 ;
        RECT 960.2000 433.6050 962.2000 435.6050 ;
        RECT 952.0500 433.6050 954.0500 435.6050 ;
        RECT 976.5000 426.5100 978.5000 428.5100 ;
        RECT 968.3500 426.5100 970.3500 428.5100 ;
        RECT 960.2000 426.5100 962.2000 428.5100 ;
        RECT 952.0500 426.5100 954.0500 428.5100 ;
        RECT 960.2000 447.7950 962.2000 449.7950 ;
        RECT 952.0500 447.7950 954.0500 449.7950 ;
        RECT 976.5000 440.7000 978.5000 442.7000 ;
        RECT 968.3500 440.7000 970.3500 442.7000 ;
        RECT 960.2000 440.7000 962.2000 442.7000 ;
        RECT 952.0500 440.7000 954.0500 442.7000 ;
        RECT 968.3500 447.7950 970.3500 449.7950 ;
        RECT 976.5000 447.7950 978.5000 449.7950 ;
        RECT 943.9000 461.9850 945.9000 463.9850 ;
        RECT 943.9000 469.0800 945.9000 471.0800 ;
        RECT 943.9000 476.1750 945.9000 478.1750 ;
        RECT 943.9000 483.2700 945.9000 485.2700 ;
        RECT 935.7500 469.0800 937.7500 471.0800 ;
        RECT 927.6000 469.0800 929.6000 471.0800 ;
        RECT 919.4500 469.0800 921.4500 471.0800 ;
        RECT 911.3000 469.0800 913.3000 471.0800 ;
        RECT 935.7500 461.9850 937.7500 463.9850 ;
        RECT 927.6000 461.9850 929.6000 463.9850 ;
        RECT 919.4500 461.9850 921.4500 463.9850 ;
        RECT 911.3000 461.9850 913.3000 463.9850 ;
        RECT 919.4500 483.2700 921.4500 485.2700 ;
        RECT 911.3000 483.2700 913.3000 485.2700 ;
        RECT 935.7500 476.1750 937.7500 478.1750 ;
        RECT 927.6000 476.1750 929.6000 478.1750 ;
        RECT 919.4500 476.1750 921.4500 478.1750 ;
        RECT 911.3000 476.1750 913.3000 478.1750 ;
        RECT 927.6000 483.2700 929.6000 485.2700 ;
        RECT 935.7500 483.2700 937.7500 485.2700 ;
        RECT 976.5000 469.0800 978.5000 471.0800 ;
        RECT 968.3500 469.0800 970.3500 471.0800 ;
        RECT 960.2000 469.0800 962.2000 471.0800 ;
        RECT 952.0500 469.0800 954.0500 471.0800 ;
        RECT 976.5000 461.9850 978.5000 463.9850 ;
        RECT 968.3500 461.9850 970.3500 463.9850 ;
        RECT 960.2000 461.9850 962.2000 463.9850 ;
        RECT 952.0500 461.9850 954.0500 463.9850 ;
        RECT 960.2000 483.2700 962.2000 485.2700 ;
        RECT 952.0500 483.2700 954.0500 485.2700 ;
        RECT 976.5000 476.1750 978.5000 478.1750 ;
        RECT 968.3500 476.1750 970.3500 478.1750 ;
        RECT 960.2000 476.1750 962.2000 478.1750 ;
        RECT 952.0500 476.1750 954.0500 478.1750 ;
        RECT 968.3500 483.2700 970.3500 485.2700 ;
        RECT 976.5000 483.2700 978.5000 485.2700 ;
        RECT 854.2500 504.5550 856.2500 506.5550 ;
        RECT 846.1000 504.5550 848.1000 506.5550 ;
        RECT 870.5500 497.4600 872.5500 499.4600 ;
        RECT 862.4000 497.4600 864.4000 499.4600 ;
        RECT 854.2500 497.4600 856.2500 499.4600 ;
        RECT 846.1000 497.4600 848.1000 499.4600 ;
        RECT 870.5500 490.3650 872.5500 492.3650 ;
        RECT 862.4000 490.3650 864.4000 492.3650 ;
        RECT 854.2500 490.3650 856.2500 492.3650 ;
        RECT 846.1000 490.3650 848.1000 492.3650 ;
        RECT 862.4000 504.5550 864.4000 506.5550 ;
        RECT 870.5500 504.5550 872.5500 506.5550 ;
        RECT 846.1000 511.6500 848.1000 513.6500 ;
        RECT 854.2500 511.6500 856.2500 513.6500 ;
        RECT 862.4000 511.6500 864.4000 513.6500 ;
        RECT 870.5500 511.6500 872.5500 513.6500 ;
        RECT 846.1000 518.7450 848.1000 520.7450 ;
        RECT 854.2500 518.7450 856.2500 520.7450 ;
        RECT 862.4000 518.7450 864.4000 520.7450 ;
        RECT 870.5500 518.7450 872.5500 520.7450 ;
        RECT 886.8500 504.5550 888.8500 506.5550 ;
        RECT 878.7000 504.5550 880.7000 506.5550 ;
        RECT 903.1500 497.4600 905.1500 499.4600 ;
        RECT 895.0000 497.4600 897.0000 499.4600 ;
        RECT 886.8500 497.4600 888.8500 499.4600 ;
        RECT 878.7000 497.4600 880.7000 499.4600 ;
        RECT 903.1500 490.3650 905.1500 492.3650 ;
        RECT 895.0000 490.3650 897.0000 492.3650 ;
        RECT 886.8500 490.3650 888.8500 492.3650 ;
        RECT 878.7000 490.3650 880.7000 492.3650 ;
        RECT 895.0000 504.5550 897.0000 506.5550 ;
        RECT 903.1500 504.5550 905.1500 506.5550 ;
        RECT 878.7000 511.6500 880.7000 513.6500 ;
        RECT 886.8500 511.6500 888.8500 513.6500 ;
        RECT 895.0000 511.6500 897.0000 513.6500 ;
        RECT 903.1500 511.6500 905.1500 513.6500 ;
        RECT 878.7000 518.7450 880.7000 520.7450 ;
        RECT 886.8500 518.7450 888.8500 520.7450 ;
        RECT 895.0000 518.7450 897.0000 520.7450 ;
        RECT 903.1500 518.7450 905.1500 520.7450 ;
        RECT 854.2500 540.0300 856.2500 542.0300 ;
        RECT 846.1000 540.0300 848.1000 542.0300 ;
        RECT 870.5500 532.9350 872.5500 534.9350 ;
        RECT 862.4000 532.9350 864.4000 534.9350 ;
        RECT 854.2500 532.9350 856.2500 534.9350 ;
        RECT 846.1000 532.9350 848.1000 534.9350 ;
        RECT 870.5500 525.8400 872.5500 527.8400 ;
        RECT 862.4000 525.8400 864.4000 527.8400 ;
        RECT 854.2500 525.8400 856.2500 527.8400 ;
        RECT 846.1000 525.8400 848.1000 527.8400 ;
        RECT 862.4000 540.0300 864.4000 542.0300 ;
        RECT 870.5500 540.0300 872.5500 542.0300 ;
        RECT 846.1000 547.1250 848.1000 549.1250 ;
        RECT 854.2500 547.1250 856.2500 549.1250 ;
        RECT 862.4000 547.1250 864.4000 549.1250 ;
        RECT 870.5500 547.1250 872.5500 549.1250 ;
        RECT 846.1000 554.2200 848.1000 556.2200 ;
        RECT 854.2500 554.2200 856.2500 556.2200 ;
        RECT 862.4000 554.2200 864.4000 556.2200 ;
        RECT 870.5500 554.2200 872.5500 556.2200 ;
        RECT 886.8500 540.0300 888.8500 542.0300 ;
        RECT 878.7000 540.0300 880.7000 542.0300 ;
        RECT 903.1500 532.9350 905.1500 534.9350 ;
        RECT 895.0000 532.9350 897.0000 534.9350 ;
        RECT 886.8500 532.9350 888.8500 534.9350 ;
        RECT 878.7000 532.9350 880.7000 534.9350 ;
        RECT 903.1500 525.8400 905.1500 527.8400 ;
        RECT 895.0000 525.8400 897.0000 527.8400 ;
        RECT 886.8500 525.8400 888.8500 527.8400 ;
        RECT 878.7000 525.8400 880.7000 527.8400 ;
        RECT 895.0000 540.0300 897.0000 542.0300 ;
        RECT 903.1500 540.0300 905.1500 542.0300 ;
        RECT 878.7000 547.1250 880.7000 549.1250 ;
        RECT 886.8500 547.1250 888.8500 549.1250 ;
        RECT 895.0000 547.1250 897.0000 549.1250 ;
        RECT 903.1500 547.1250 905.1500 549.1250 ;
        RECT 878.7000 554.2200 880.7000 556.2200 ;
        RECT 886.8500 554.2200 888.8500 556.2200 ;
        RECT 895.0000 554.2200 897.0000 556.2200 ;
        RECT 903.1500 554.2200 905.1500 556.2200 ;
        RECT 943.9000 490.3650 945.9000 492.3650 ;
        RECT 943.9000 497.4600 945.9000 499.4600 ;
        RECT 943.9000 504.5550 945.9000 506.5550 ;
        RECT 943.9000 511.6500 945.9000 513.6500 ;
        RECT 943.9000 518.7450 945.9000 520.7450 ;
        RECT 919.4500 504.5550 921.4500 506.5550 ;
        RECT 911.3000 504.5550 913.3000 506.5550 ;
        RECT 935.7500 497.4600 937.7500 499.4600 ;
        RECT 927.6000 497.4600 929.6000 499.4600 ;
        RECT 919.4500 497.4600 921.4500 499.4600 ;
        RECT 911.3000 497.4600 913.3000 499.4600 ;
        RECT 935.7500 490.3650 937.7500 492.3650 ;
        RECT 927.6000 490.3650 929.6000 492.3650 ;
        RECT 919.4500 490.3650 921.4500 492.3650 ;
        RECT 911.3000 490.3650 913.3000 492.3650 ;
        RECT 927.6000 504.5550 929.6000 506.5550 ;
        RECT 935.7500 504.5550 937.7500 506.5550 ;
        RECT 911.3000 511.6500 913.3000 513.6500 ;
        RECT 919.4500 511.6500 921.4500 513.6500 ;
        RECT 927.6000 511.6500 929.6000 513.6500 ;
        RECT 935.7500 511.6500 937.7500 513.6500 ;
        RECT 911.3000 518.7450 913.3000 520.7450 ;
        RECT 919.4500 518.7450 921.4500 520.7450 ;
        RECT 927.6000 518.7450 929.6000 520.7450 ;
        RECT 935.7500 518.7450 937.7500 520.7450 ;
        RECT 960.2000 504.5550 962.2000 506.5550 ;
        RECT 952.0500 504.5550 954.0500 506.5550 ;
        RECT 976.5000 497.4600 978.5000 499.4600 ;
        RECT 968.3500 497.4600 970.3500 499.4600 ;
        RECT 960.2000 497.4600 962.2000 499.4600 ;
        RECT 952.0500 497.4600 954.0500 499.4600 ;
        RECT 976.5000 490.3650 978.5000 492.3650 ;
        RECT 968.3500 490.3650 970.3500 492.3650 ;
        RECT 960.2000 490.3650 962.2000 492.3650 ;
        RECT 952.0500 490.3650 954.0500 492.3650 ;
        RECT 968.3500 504.5550 970.3500 506.5550 ;
        RECT 976.5000 504.5550 978.5000 506.5550 ;
        RECT 952.0500 511.6500 954.0500 513.6500 ;
        RECT 960.2000 511.6500 962.2000 513.6500 ;
        RECT 968.3500 511.6500 970.3500 513.6500 ;
        RECT 976.5000 511.6500 978.5000 513.6500 ;
        RECT 952.0500 518.7450 954.0500 520.7450 ;
        RECT 960.2000 518.7450 962.2000 520.7450 ;
        RECT 968.3500 518.7450 970.3500 520.7450 ;
        RECT 976.5000 518.7450 978.5000 520.7450 ;
        RECT 943.9000 525.8400 945.9000 527.8400 ;
        RECT 943.9000 532.9350 945.9000 534.9350 ;
        RECT 943.9000 540.0300 945.9000 542.0300 ;
        RECT 943.9000 547.1250 945.9000 549.1250 ;
        RECT 943.9000 554.2200 945.9000 556.2200 ;
        RECT 919.4500 540.0300 921.4500 542.0300 ;
        RECT 911.3000 540.0300 913.3000 542.0300 ;
        RECT 935.7500 532.9350 937.7500 534.9350 ;
        RECT 927.6000 532.9350 929.6000 534.9350 ;
        RECT 919.4500 532.9350 921.4500 534.9350 ;
        RECT 911.3000 532.9350 913.3000 534.9350 ;
        RECT 935.7500 525.8400 937.7500 527.8400 ;
        RECT 927.6000 525.8400 929.6000 527.8400 ;
        RECT 919.4500 525.8400 921.4500 527.8400 ;
        RECT 911.3000 525.8400 913.3000 527.8400 ;
        RECT 927.6000 540.0300 929.6000 542.0300 ;
        RECT 935.7500 540.0300 937.7500 542.0300 ;
        RECT 911.3000 547.1250 913.3000 549.1250 ;
        RECT 919.4500 547.1250 921.4500 549.1250 ;
        RECT 927.6000 547.1250 929.6000 549.1250 ;
        RECT 935.7500 547.1250 937.7500 549.1250 ;
        RECT 911.3000 554.2200 913.3000 556.2200 ;
        RECT 919.4500 554.2200 921.4500 556.2200 ;
        RECT 927.6000 554.2200 929.6000 556.2200 ;
        RECT 935.7500 554.2200 937.7500 556.2200 ;
        RECT 960.2000 540.0300 962.2000 542.0300 ;
        RECT 952.0500 540.0300 954.0500 542.0300 ;
        RECT 976.5000 532.9350 978.5000 534.9350 ;
        RECT 968.3500 532.9350 970.3500 534.9350 ;
        RECT 960.2000 532.9350 962.2000 534.9350 ;
        RECT 952.0500 532.9350 954.0500 534.9350 ;
        RECT 976.5000 525.8400 978.5000 527.8400 ;
        RECT 968.3500 525.8400 970.3500 527.8400 ;
        RECT 960.2000 525.8400 962.2000 527.8400 ;
        RECT 952.0500 525.8400 954.0500 527.8400 ;
        RECT 968.3500 540.0300 970.3500 542.0300 ;
        RECT 976.5000 540.0300 978.5000 542.0300 ;
        RECT 952.0500 547.1250 954.0500 549.1250 ;
        RECT 960.2000 547.1250 962.2000 549.1250 ;
        RECT 968.3500 547.1250 970.3500 549.1250 ;
        RECT 976.5000 547.1250 978.5000 549.1250 ;
        RECT 952.0500 554.2200 954.0500 556.2200 ;
        RECT 960.2000 554.2200 962.2000 556.2200 ;
        RECT 968.3500 554.2200 970.3500 556.2200 ;
        RECT 976.5000 554.2200 978.5000 556.2200 ;
        RECT 1049.8500 426.5100 1051.8500 428.5100 ;
        RECT 1049.8500 433.6050 1051.8500 435.6050 ;
        RECT 1049.8500 440.7000 1051.8500 442.7000 ;
        RECT 1049.8500 447.7950 1051.8500 449.7950 ;
        RECT 1049.8500 454.8900 1051.8500 456.8900 ;
        RECT 1049.8500 461.9850 1051.8500 463.9850 ;
        RECT 1049.8500 469.0800 1051.8500 471.0800 ;
        RECT 1049.8500 476.1750 1051.8500 478.1750 ;
        RECT 1049.8500 483.2700 1051.8500 485.2700 ;
        RECT 984.6500 454.8900 986.6500 456.8900 ;
        RECT 992.8000 454.8900 994.8000 456.8900 ;
        RECT 1000.9500 454.8900 1002.9500 456.8900 ;
        RECT 1009.1000 454.8900 1011.1000 456.8900 ;
        RECT 1017.2500 454.8900 1019.2500 456.8900 ;
        RECT 1025.4000 454.8900 1027.4000 456.8900 ;
        RECT 1033.5500 454.8900 1035.5500 456.8900 ;
        RECT 1041.7000 454.8900 1043.7000 456.8900 ;
        RECT 1009.1000 433.6050 1011.1000 435.6050 ;
        RECT 1000.9500 433.6050 1002.9500 435.6050 ;
        RECT 992.8000 433.6050 994.8000 435.6050 ;
        RECT 984.6500 433.6050 986.6500 435.6050 ;
        RECT 1009.1000 426.5100 1011.1000 428.5100 ;
        RECT 1000.9500 426.5100 1002.9500 428.5100 ;
        RECT 992.8000 426.5100 994.8000 428.5100 ;
        RECT 984.6500 426.5100 986.6500 428.5100 ;
        RECT 992.8000 447.7950 994.8000 449.7950 ;
        RECT 984.6500 447.7950 986.6500 449.7950 ;
        RECT 1009.1000 440.7000 1011.1000 442.7000 ;
        RECT 1000.9500 440.7000 1002.9500 442.7000 ;
        RECT 992.8000 440.7000 994.8000 442.7000 ;
        RECT 984.6500 440.7000 986.6500 442.7000 ;
        RECT 1000.9500 447.7950 1002.9500 449.7950 ;
        RECT 1009.1000 447.7950 1011.1000 449.7950 ;
        RECT 1041.7000 433.6050 1043.7000 435.6050 ;
        RECT 1033.5500 433.6050 1035.5500 435.6050 ;
        RECT 1025.4000 433.6050 1027.4000 435.6050 ;
        RECT 1017.2500 433.6050 1019.2500 435.6050 ;
        RECT 1041.7000 426.5100 1043.7000 428.5100 ;
        RECT 1033.5500 426.5100 1035.5500 428.5100 ;
        RECT 1025.4000 426.5100 1027.4000 428.5100 ;
        RECT 1017.2500 426.5100 1019.2500 428.5100 ;
        RECT 1025.4000 447.7950 1027.4000 449.7950 ;
        RECT 1017.2500 447.7950 1019.2500 449.7950 ;
        RECT 1041.7000 440.7000 1043.7000 442.7000 ;
        RECT 1033.5500 440.7000 1035.5500 442.7000 ;
        RECT 1025.4000 440.7000 1027.4000 442.7000 ;
        RECT 1017.2500 440.7000 1019.2500 442.7000 ;
        RECT 1033.5500 447.7950 1035.5500 449.7950 ;
        RECT 1041.7000 447.7950 1043.7000 449.7950 ;
        RECT 1009.1000 469.0800 1011.1000 471.0800 ;
        RECT 1000.9500 469.0800 1002.9500 471.0800 ;
        RECT 992.8000 469.0800 994.8000 471.0800 ;
        RECT 984.6500 469.0800 986.6500 471.0800 ;
        RECT 1009.1000 461.9850 1011.1000 463.9850 ;
        RECT 1000.9500 461.9850 1002.9500 463.9850 ;
        RECT 992.8000 461.9850 994.8000 463.9850 ;
        RECT 984.6500 461.9850 986.6500 463.9850 ;
        RECT 992.8000 483.2700 994.8000 485.2700 ;
        RECT 984.6500 483.2700 986.6500 485.2700 ;
        RECT 1009.1000 476.1750 1011.1000 478.1750 ;
        RECT 1000.9500 476.1750 1002.9500 478.1750 ;
        RECT 992.8000 476.1750 994.8000 478.1750 ;
        RECT 984.6500 476.1750 986.6500 478.1750 ;
        RECT 1000.9500 483.2700 1002.9500 485.2700 ;
        RECT 1009.1000 483.2700 1011.1000 485.2700 ;
        RECT 1041.7000 469.0800 1043.7000 471.0800 ;
        RECT 1033.5500 469.0800 1035.5500 471.0800 ;
        RECT 1025.4000 469.0800 1027.4000 471.0800 ;
        RECT 1017.2500 469.0800 1019.2500 471.0800 ;
        RECT 1041.7000 461.9850 1043.7000 463.9850 ;
        RECT 1033.5500 461.9850 1035.5500 463.9850 ;
        RECT 1025.4000 461.9850 1027.4000 463.9850 ;
        RECT 1017.2500 461.9850 1019.2500 463.9850 ;
        RECT 1025.4000 483.2700 1027.4000 485.2700 ;
        RECT 1017.2500 483.2700 1019.2500 485.2700 ;
        RECT 1041.7000 476.1750 1043.7000 478.1750 ;
        RECT 1033.5500 476.1750 1035.5500 478.1750 ;
        RECT 1025.4000 476.1750 1027.4000 478.1750 ;
        RECT 1017.2500 476.1750 1019.2500 478.1750 ;
        RECT 1033.5500 483.2700 1035.5500 485.2700 ;
        RECT 1041.7000 483.2700 1043.7000 485.2700 ;
        RECT 1074.0000 454.8900 1076.0000 456.8900 ;
        RECT 1112.0000 454.8900 1114.0000 456.8900 ;
        RECT 1058.0000 454.8900 1060.0000 456.8900 ;
        RECT 1058.0000 433.6050 1060.0000 435.6050 ;
        RECT 1058.0000 426.5100 1060.0000 428.5100 ;
        RECT 1074.0000 426.5100 1076.0000 428.5100 ;
        RECT 1074.0000 433.6050 1076.0000 435.6050 ;
        RECT 1058.0000 447.7950 1060.0000 449.7950 ;
        RECT 1058.0000 440.7000 1060.0000 442.7000 ;
        RECT 1074.0000 440.7000 1076.0000 442.7000 ;
        RECT 1074.0000 447.7950 1076.0000 449.7950 ;
        RECT 1112.0000 426.5100 1114.0000 428.5100 ;
        RECT 1112.0000 433.6050 1114.0000 435.6050 ;
        RECT 1112.0000 440.7000 1114.0000 442.7000 ;
        RECT 1112.0000 447.7950 1114.0000 449.7950 ;
        RECT 1058.0000 469.0800 1060.0000 471.0800 ;
        RECT 1058.0000 461.9850 1060.0000 463.9850 ;
        RECT 1074.0000 469.0800 1076.0000 471.0800 ;
        RECT 1074.0000 461.9850 1076.0000 463.9850 ;
        RECT 1058.0000 483.2700 1060.0000 485.2700 ;
        RECT 1058.0000 476.1750 1060.0000 478.1750 ;
        RECT 1074.0000 483.2700 1076.0000 485.2700 ;
        RECT 1074.0000 476.1750 1076.0000 478.1750 ;
        RECT 1112.0000 461.9850 1114.0000 463.9850 ;
        RECT 1112.0000 469.0800 1114.0000 471.0800 ;
        RECT 1112.0000 476.1750 1114.0000 478.1750 ;
        RECT 1112.0000 483.2700 1114.0000 485.2700 ;
        RECT 1049.8500 490.3650 1051.8500 492.3650 ;
        RECT 1049.8500 497.4600 1051.8500 499.4600 ;
        RECT 1049.8500 504.5550 1051.8500 506.5550 ;
        RECT 1049.8500 511.6500 1051.8500 513.6500 ;
        RECT 1049.8500 518.7450 1051.8500 520.7450 ;
        RECT 1049.8500 525.8400 1051.8500 527.8400 ;
        RECT 1049.8500 532.9350 1051.8500 534.9350 ;
        RECT 1049.8500 540.0300 1051.8500 542.0300 ;
        RECT 1049.8500 547.1250 1051.8500 549.1250 ;
        RECT 1049.8500 554.2200 1051.8500 556.2200 ;
        RECT 992.8000 504.5550 994.8000 506.5550 ;
        RECT 984.6500 504.5550 986.6500 506.5550 ;
        RECT 1009.1000 497.4600 1011.1000 499.4600 ;
        RECT 1000.9500 497.4600 1002.9500 499.4600 ;
        RECT 992.8000 497.4600 994.8000 499.4600 ;
        RECT 984.6500 497.4600 986.6500 499.4600 ;
        RECT 1009.1000 490.3650 1011.1000 492.3650 ;
        RECT 1000.9500 490.3650 1002.9500 492.3650 ;
        RECT 992.8000 490.3650 994.8000 492.3650 ;
        RECT 984.6500 490.3650 986.6500 492.3650 ;
        RECT 1000.9500 504.5550 1002.9500 506.5550 ;
        RECT 1009.1000 504.5550 1011.1000 506.5550 ;
        RECT 984.6500 511.6500 986.6500 513.6500 ;
        RECT 992.8000 511.6500 994.8000 513.6500 ;
        RECT 1000.9500 511.6500 1002.9500 513.6500 ;
        RECT 1009.1000 511.6500 1011.1000 513.6500 ;
        RECT 984.6500 518.7450 986.6500 520.7450 ;
        RECT 992.8000 518.7450 994.8000 520.7450 ;
        RECT 1000.9500 518.7450 1002.9500 520.7450 ;
        RECT 1009.1000 518.7450 1011.1000 520.7450 ;
        RECT 1025.4000 504.5550 1027.4000 506.5550 ;
        RECT 1017.2500 504.5550 1019.2500 506.5550 ;
        RECT 1041.7000 497.4600 1043.7000 499.4600 ;
        RECT 1033.5500 497.4600 1035.5500 499.4600 ;
        RECT 1025.4000 497.4600 1027.4000 499.4600 ;
        RECT 1017.2500 497.4600 1019.2500 499.4600 ;
        RECT 1041.7000 490.3650 1043.7000 492.3650 ;
        RECT 1033.5500 490.3650 1035.5500 492.3650 ;
        RECT 1025.4000 490.3650 1027.4000 492.3650 ;
        RECT 1017.2500 490.3650 1019.2500 492.3650 ;
        RECT 1033.5500 504.5550 1035.5500 506.5550 ;
        RECT 1041.7000 504.5550 1043.7000 506.5550 ;
        RECT 1017.2500 511.6500 1019.2500 513.6500 ;
        RECT 1025.4000 511.6500 1027.4000 513.6500 ;
        RECT 1033.5500 511.6500 1035.5500 513.6500 ;
        RECT 1041.7000 511.6500 1043.7000 513.6500 ;
        RECT 1017.2500 518.7450 1019.2500 520.7450 ;
        RECT 1025.4000 518.7450 1027.4000 520.7450 ;
        RECT 1033.5500 518.7450 1035.5500 520.7450 ;
        RECT 1041.7000 518.7450 1043.7000 520.7450 ;
        RECT 992.8000 540.0300 994.8000 542.0300 ;
        RECT 984.6500 540.0300 986.6500 542.0300 ;
        RECT 1009.1000 532.9350 1011.1000 534.9350 ;
        RECT 1000.9500 532.9350 1002.9500 534.9350 ;
        RECT 992.8000 532.9350 994.8000 534.9350 ;
        RECT 984.6500 532.9350 986.6500 534.9350 ;
        RECT 1009.1000 525.8400 1011.1000 527.8400 ;
        RECT 1000.9500 525.8400 1002.9500 527.8400 ;
        RECT 992.8000 525.8400 994.8000 527.8400 ;
        RECT 984.6500 525.8400 986.6500 527.8400 ;
        RECT 1000.9500 540.0300 1002.9500 542.0300 ;
        RECT 1009.1000 540.0300 1011.1000 542.0300 ;
        RECT 984.6500 547.1250 986.6500 549.1250 ;
        RECT 992.8000 547.1250 994.8000 549.1250 ;
        RECT 1000.9500 547.1250 1002.9500 549.1250 ;
        RECT 1009.1000 547.1250 1011.1000 549.1250 ;
        RECT 984.6500 554.2200 986.6500 556.2200 ;
        RECT 992.8000 554.2200 994.8000 556.2200 ;
        RECT 1000.9500 554.2200 1002.9500 556.2200 ;
        RECT 1009.1000 554.2200 1011.1000 556.2200 ;
        RECT 1025.4000 540.0300 1027.4000 542.0300 ;
        RECT 1017.2500 540.0300 1019.2500 542.0300 ;
        RECT 1041.7000 532.9350 1043.7000 534.9350 ;
        RECT 1033.5500 532.9350 1035.5500 534.9350 ;
        RECT 1025.4000 532.9350 1027.4000 534.9350 ;
        RECT 1017.2500 532.9350 1019.2500 534.9350 ;
        RECT 1041.7000 525.8400 1043.7000 527.8400 ;
        RECT 1033.5500 525.8400 1035.5500 527.8400 ;
        RECT 1025.4000 525.8400 1027.4000 527.8400 ;
        RECT 1017.2500 525.8400 1019.2500 527.8400 ;
        RECT 1033.5500 540.0300 1035.5500 542.0300 ;
        RECT 1041.7000 540.0300 1043.7000 542.0300 ;
        RECT 1017.2500 547.1250 1019.2500 549.1250 ;
        RECT 1025.4000 547.1250 1027.4000 549.1250 ;
        RECT 1033.5500 547.1250 1035.5500 549.1250 ;
        RECT 1041.7000 547.1250 1043.7000 549.1250 ;
        RECT 1017.2500 554.2200 1019.2500 556.2200 ;
        RECT 1025.4000 554.2200 1027.4000 556.2200 ;
        RECT 1033.5500 554.2200 1035.5500 556.2200 ;
        RECT 1041.7000 554.2200 1043.7000 556.2200 ;
        RECT 1058.0000 490.3650 1060.0000 492.3650 ;
        RECT 1058.0000 497.4600 1060.0000 499.4600 ;
        RECT 1058.0000 504.5550 1060.0000 506.5550 ;
        RECT 1074.0000 497.4600 1076.0000 499.4600 ;
        RECT 1074.0000 490.3650 1076.0000 492.3650 ;
        RECT 1074.0000 504.5550 1076.0000 506.5550 ;
        RECT 1058.0000 518.7450 1060.0000 520.7450 ;
        RECT 1058.0000 511.6500 1060.0000 513.6500 ;
        RECT 1074.0000 511.6500 1076.0000 513.6500 ;
        RECT 1074.0000 518.7450 1076.0000 520.7450 ;
        RECT 1112.0000 497.4600 1114.0000 499.4600 ;
        RECT 1112.0000 490.3650 1114.0000 492.3650 ;
        RECT 1112.0000 504.5550 1114.0000 506.5550 ;
        RECT 1112.0000 511.6500 1114.0000 513.6500 ;
        RECT 1112.0000 518.7450 1114.0000 520.7450 ;
        RECT 1058.0000 532.9350 1060.0000 534.9350 ;
        RECT 1058.0000 525.8400 1060.0000 527.8400 ;
        RECT 1058.0000 540.0300 1060.0000 542.0300 ;
        RECT 1074.0000 532.9350 1076.0000 534.9350 ;
        RECT 1074.0000 525.8400 1076.0000 527.8400 ;
        RECT 1074.0000 540.0300 1076.0000 542.0300 ;
        RECT 1058.0000 554.2200 1060.0000 556.2200 ;
        RECT 1058.0000 547.1250 1060.0000 549.1250 ;
        RECT 1074.0000 547.1250 1076.0000 549.1250 ;
        RECT 1074.0000 554.2200 1076.0000 556.2200 ;
        RECT 1112.0000 532.9350 1114.0000 534.9350 ;
        RECT 1112.0000 525.8400 1114.0000 527.8400 ;
        RECT 1112.0000 540.0300 1114.0000 542.0300 ;
        RECT 1112.0000 547.1250 1114.0000 549.1250 ;
        RECT 1112.0000 554.2200 1114.0000 556.2200 ;
        RECT 6.0000 838.0200 8.0000 840.0200 ;
        RECT 68.5150 561.3150 70.5150 563.3150 ;
        RECT 68.5150 568.4100 70.5150 570.4100 ;
        RECT 68.5150 575.5050 70.5150 577.5050 ;
        RECT 68.5150 582.6000 70.5150 584.6000 ;
        RECT 68.5150 589.6950 70.5150 591.6950 ;
        RECT 68.5150 596.7900 70.5150 598.7900 ;
        RECT 68.5150 603.8850 70.5150 605.8850 ;
        RECT 68.5150 610.9800 70.5150 612.9800 ;
        RECT 68.5150 618.0750 70.5150 620.0750 ;
        RECT 68.5150 625.1700 70.5150 627.1700 ;
        RECT 6.0000 575.5050 8.0000 577.5050 ;
        RECT 6.0000 568.4100 8.0000 570.4100 ;
        RECT 6.0000 561.3150 8.0000 563.3150 ;
        RECT 6.0000 582.6000 8.0000 584.6000 ;
        RECT 6.0000 589.6950 8.0000 591.6950 ;
        RECT 44.0000 575.5050 46.0000 577.5050 ;
        RECT 60.0000 575.5050 62.0000 577.5050 ;
        RECT 44.0000 561.3150 46.0000 563.3150 ;
        RECT 44.0000 568.4100 46.0000 570.4100 ;
        RECT 60.0000 568.4100 62.0000 570.4100 ;
        RECT 60.0000 561.3150 62.0000 563.3150 ;
        RECT 44.0000 589.6950 46.0000 591.6950 ;
        RECT 44.0000 582.6000 46.0000 584.6000 ;
        RECT 60.0000 582.6000 62.0000 584.6000 ;
        RECT 60.0000 589.6950 62.0000 591.6950 ;
        RECT 6.0000 610.9800 8.0000 612.9800 ;
        RECT 6.0000 596.7900 8.0000 598.7900 ;
        RECT 6.0000 603.8850 8.0000 605.8850 ;
        RECT 6.0000 618.0750 8.0000 620.0750 ;
        RECT 6.0000 625.1700 8.0000 627.1700 ;
        RECT 44.0000 610.9800 46.0000 612.9800 ;
        RECT 60.0000 610.9800 62.0000 612.9800 ;
        RECT 44.0000 603.8850 46.0000 605.8850 ;
        RECT 44.0000 596.7900 46.0000 598.7900 ;
        RECT 60.0000 596.7900 62.0000 598.7900 ;
        RECT 60.0000 603.8850 62.0000 605.8850 ;
        RECT 44.0000 618.0750 46.0000 620.0750 ;
        RECT 44.0000 625.1700 46.0000 627.1700 ;
        RECT 60.0000 625.1700 62.0000 627.1700 ;
        RECT 60.0000 618.0750 62.0000 620.0750 ;
        RECT 77.0300 575.5050 79.0300 577.5050 ;
        RECT 85.5450 575.5050 87.5450 577.5050 ;
        RECT 94.0600 575.5050 96.0600 577.5050 ;
        RECT 102.5750 575.5050 104.5750 577.5050 ;
        RECT 102.5750 568.4100 104.5750 570.4100 ;
        RECT 94.0600 568.4100 96.0600 570.4100 ;
        RECT 85.5450 568.4100 87.5450 570.4100 ;
        RECT 77.0300 568.4100 79.0300 570.4100 ;
        RECT 102.5750 561.3150 104.5750 563.3150 ;
        RECT 94.0600 561.3150 96.0600 563.3150 ;
        RECT 85.5450 561.3150 87.5450 563.3150 ;
        RECT 77.0300 561.3150 79.0300 563.3150 ;
        RECT 77.0300 582.6000 79.0300 584.6000 ;
        RECT 85.5450 582.6000 87.5450 584.6000 ;
        RECT 94.0600 582.6000 96.0600 584.6000 ;
        RECT 102.5750 582.6000 104.5750 584.6000 ;
        RECT 77.0300 589.6950 79.0300 591.6950 ;
        RECT 85.5450 589.6950 87.5450 591.6950 ;
        RECT 94.0600 589.6950 96.0600 591.6950 ;
        RECT 102.5750 589.6950 104.5750 591.6950 ;
        RECT 111.0900 575.5050 113.0900 577.5050 ;
        RECT 119.6050 575.5050 121.6050 577.5050 ;
        RECT 128.1200 575.5050 130.1200 577.5050 ;
        RECT 136.6350 575.5050 138.6350 577.5050 ;
        RECT 136.6350 568.4100 138.6350 570.4100 ;
        RECT 128.1200 568.4100 130.1200 570.4100 ;
        RECT 119.6050 568.4100 121.6050 570.4100 ;
        RECT 111.0900 568.4100 113.0900 570.4100 ;
        RECT 136.6350 561.3150 138.6350 563.3150 ;
        RECT 128.1200 561.3150 130.1200 563.3150 ;
        RECT 119.6050 561.3150 121.6050 563.3150 ;
        RECT 111.0900 561.3150 113.0900 563.3150 ;
        RECT 111.0900 582.6000 113.0900 584.6000 ;
        RECT 119.6050 582.6000 121.6050 584.6000 ;
        RECT 128.1200 582.6000 130.1200 584.6000 ;
        RECT 136.6350 582.6000 138.6350 584.6000 ;
        RECT 111.0900 589.6950 113.0900 591.6950 ;
        RECT 119.6050 589.6950 121.6050 591.6950 ;
        RECT 128.1200 589.6950 130.1200 591.6950 ;
        RECT 136.6350 589.6950 138.6350 591.6950 ;
        RECT 77.0300 610.9800 79.0300 612.9800 ;
        RECT 85.5450 610.9800 87.5450 612.9800 ;
        RECT 94.0600 610.9800 96.0600 612.9800 ;
        RECT 102.5750 610.9800 104.5750 612.9800 ;
        RECT 102.5750 603.8850 104.5750 605.8850 ;
        RECT 94.0600 603.8850 96.0600 605.8850 ;
        RECT 85.5450 603.8850 87.5450 605.8850 ;
        RECT 77.0300 603.8850 79.0300 605.8850 ;
        RECT 102.5750 596.7900 104.5750 598.7900 ;
        RECT 94.0600 596.7900 96.0600 598.7900 ;
        RECT 85.5450 596.7900 87.5450 598.7900 ;
        RECT 77.0300 596.7900 79.0300 598.7900 ;
        RECT 77.0300 618.0750 79.0300 620.0750 ;
        RECT 85.5450 618.0750 87.5450 620.0750 ;
        RECT 94.0600 618.0750 96.0600 620.0750 ;
        RECT 102.5750 618.0750 104.5750 620.0750 ;
        RECT 77.0300 625.1700 79.0300 627.1700 ;
        RECT 85.5450 625.1700 87.5450 627.1700 ;
        RECT 94.0600 625.1700 96.0600 627.1700 ;
        RECT 102.5750 625.1700 104.5750 627.1700 ;
        RECT 111.0900 610.9800 113.0900 612.9800 ;
        RECT 119.6050 610.9800 121.6050 612.9800 ;
        RECT 128.1200 610.9800 130.1200 612.9800 ;
        RECT 136.6350 610.9800 138.6350 612.9800 ;
        RECT 136.6350 603.8850 138.6350 605.8850 ;
        RECT 128.1200 603.8850 130.1200 605.8850 ;
        RECT 119.6050 603.8850 121.6050 605.8850 ;
        RECT 111.0900 603.8850 113.0900 605.8850 ;
        RECT 136.6350 596.7900 138.6350 598.7900 ;
        RECT 128.1200 596.7900 130.1200 598.7900 ;
        RECT 119.6050 596.7900 121.6050 598.7900 ;
        RECT 111.0900 596.7900 113.0900 598.7900 ;
        RECT 111.0900 618.0750 113.0900 620.0750 ;
        RECT 119.6050 618.0750 121.6050 620.0750 ;
        RECT 128.1200 618.0750 130.1200 620.0750 ;
        RECT 136.6350 618.0750 138.6350 620.0750 ;
        RECT 111.0900 625.1700 113.0900 627.1700 ;
        RECT 119.6050 625.1700 121.6050 627.1700 ;
        RECT 128.1200 625.1700 130.1200 627.1700 ;
        RECT 136.6350 625.1700 138.6350 627.1700 ;
        RECT 68.5150 632.2650 70.5150 634.2650 ;
        RECT 68.5150 639.3600 70.5150 641.3600 ;
        RECT 68.5150 646.4550 70.5150 648.4550 ;
        RECT 68.5150 653.5500 70.5150 655.5500 ;
        RECT 68.5150 660.6450 70.5150 662.6450 ;
        RECT 68.5150 667.7400 70.5150 669.7400 ;
        RECT 68.5150 674.8350 70.5150 676.8350 ;
        RECT 6.0000 646.4550 8.0000 648.4550 ;
        RECT 6.0000 632.2650 8.0000 634.2650 ;
        RECT 6.0000 639.3600 8.0000 641.3600 ;
        RECT 6.0000 660.6450 8.0000 662.6450 ;
        RECT 6.0000 653.5500 8.0000 655.5500 ;
        RECT 44.0000 646.4550 46.0000 648.4550 ;
        RECT 60.0000 646.4550 62.0000 648.4550 ;
        RECT 44.0000 632.2650 46.0000 634.2650 ;
        RECT 44.0000 639.3600 46.0000 641.3600 ;
        RECT 60.0000 639.3600 62.0000 641.3600 ;
        RECT 60.0000 632.2650 62.0000 634.2650 ;
        RECT 44.0000 660.6450 46.0000 662.6450 ;
        RECT 44.0000 653.5500 46.0000 655.5500 ;
        RECT 60.0000 653.5500 62.0000 655.5500 ;
        RECT 60.0000 660.6450 62.0000 662.6450 ;
        RECT 6.0000 681.9300 8.0000 683.9300 ;
        RECT 6.0000 667.7400 8.0000 669.7400 ;
        RECT 6.0000 674.8350 8.0000 676.8350 ;
        RECT 6.0000 689.0250 8.0000 691.0250 ;
        RECT 6.0000 696.1200 8.0000 698.1200 ;
        RECT 44.0000 681.9300 46.0000 683.9300 ;
        RECT 44.0000 667.7400 46.0000 669.7400 ;
        RECT 44.0000 674.8350 46.0000 676.8350 ;
        RECT 60.0000 674.8350 62.0000 676.8350 ;
        RECT 60.0000 667.7400 62.0000 669.7400 ;
        RECT 60.0000 678.0000 62.0000 680.0000 ;
        RECT 44.0000 689.0250 46.0000 691.0250 ;
        RECT 77.0300 646.4550 79.0300 648.4550 ;
        RECT 85.5450 646.4550 87.5450 648.4550 ;
        RECT 94.0600 646.4550 96.0600 648.4550 ;
        RECT 102.5750 646.4550 104.5750 648.4550 ;
        RECT 102.5750 639.3600 104.5750 641.3600 ;
        RECT 94.0600 639.3600 96.0600 641.3600 ;
        RECT 85.5450 639.3600 87.5450 641.3600 ;
        RECT 77.0300 639.3600 79.0300 641.3600 ;
        RECT 102.5750 632.2650 104.5750 634.2650 ;
        RECT 94.0600 632.2650 96.0600 634.2650 ;
        RECT 85.5450 632.2650 87.5450 634.2650 ;
        RECT 77.0300 632.2650 79.0300 634.2650 ;
        RECT 77.0300 653.5500 79.0300 655.5500 ;
        RECT 85.5450 653.5500 87.5450 655.5500 ;
        RECT 94.0600 653.5500 96.0600 655.5500 ;
        RECT 102.5750 653.5500 104.5750 655.5500 ;
        RECT 77.0300 660.6450 79.0300 662.6450 ;
        RECT 85.5450 660.6450 87.5450 662.6450 ;
        RECT 94.0600 660.6450 96.0600 662.6450 ;
        RECT 102.5750 660.6450 104.5750 662.6450 ;
        RECT 111.0900 646.4550 113.0900 648.4550 ;
        RECT 119.6050 646.4550 121.6050 648.4550 ;
        RECT 128.1200 646.4550 130.1200 648.4550 ;
        RECT 136.6350 646.4550 138.6350 648.4550 ;
        RECT 136.6350 639.3600 138.6350 641.3600 ;
        RECT 128.1200 639.3600 130.1200 641.3600 ;
        RECT 119.6050 639.3600 121.6050 641.3600 ;
        RECT 111.0900 639.3600 113.0900 641.3600 ;
        RECT 136.6350 632.2650 138.6350 634.2650 ;
        RECT 128.1200 632.2650 130.1200 634.2650 ;
        RECT 119.6050 632.2650 121.6050 634.2650 ;
        RECT 111.0900 632.2650 113.0900 634.2650 ;
        RECT 111.0900 653.5500 113.0900 655.5500 ;
        RECT 119.6050 653.5500 121.6050 655.5500 ;
        RECT 128.1200 653.5500 130.1200 655.5500 ;
        RECT 136.6350 653.5500 138.6350 655.5500 ;
        RECT 111.0900 660.6450 113.0900 662.6450 ;
        RECT 119.6050 660.6450 121.6050 662.6450 ;
        RECT 128.1200 660.6450 130.1200 662.6450 ;
        RECT 136.6350 660.6450 138.6350 662.6450 ;
        RECT 102.5750 674.8350 104.5750 676.8350 ;
        RECT 94.0600 674.8350 96.0600 676.8350 ;
        RECT 85.5450 674.8350 87.5450 676.8350 ;
        RECT 77.0300 674.8350 79.0300 676.8350 ;
        RECT 102.5750 667.7400 104.5750 669.7400 ;
        RECT 94.0600 667.7400 96.0600 669.7400 ;
        RECT 85.5450 667.7400 87.5450 669.7400 ;
        RECT 77.0300 667.7400 79.0300 669.7400 ;
        RECT 119.6050 674.8350 121.6050 676.8350 ;
        RECT 111.0900 674.8350 113.0900 676.8350 ;
        RECT 136.6350 667.7400 138.6350 669.7400 ;
        RECT 128.1200 667.7400 130.1200 669.7400 ;
        RECT 119.6050 667.7400 121.6050 669.7400 ;
        RECT 111.0900 667.7400 113.0900 669.7400 ;
        RECT 128.1200 674.8350 130.1200 676.8350 ;
        RECT 136.6350 674.8350 138.6350 676.8350 ;
        RECT 145.1500 575.5050 147.1500 577.5050 ;
        RECT 153.6650 575.5050 155.6650 577.5050 ;
        RECT 162.1800 575.5050 164.1800 577.5050 ;
        RECT 170.6950 575.5050 172.6950 577.5050 ;
        RECT 170.6950 568.4100 172.6950 570.4100 ;
        RECT 162.1800 568.4100 164.1800 570.4100 ;
        RECT 153.6650 568.4100 155.6650 570.4100 ;
        RECT 145.1500 568.4100 147.1500 570.4100 ;
        RECT 170.6950 561.3150 172.6950 563.3150 ;
        RECT 162.1800 561.3150 164.1800 563.3150 ;
        RECT 153.6650 561.3150 155.6650 563.3150 ;
        RECT 145.1500 561.3150 147.1500 563.3150 ;
        RECT 145.1500 582.6000 147.1500 584.6000 ;
        RECT 153.6650 582.6000 155.6650 584.6000 ;
        RECT 162.1800 582.6000 164.1800 584.6000 ;
        RECT 170.6950 582.6000 172.6950 584.6000 ;
        RECT 145.1500 589.6950 147.1500 591.6950 ;
        RECT 153.6650 589.6950 155.6650 591.6950 ;
        RECT 162.1800 589.6950 164.1800 591.6950 ;
        RECT 170.6950 589.6950 172.6950 591.6950 ;
        RECT 179.2100 575.5050 181.2100 577.5050 ;
        RECT 187.7250 575.5050 189.7250 577.5050 ;
        RECT 196.2400 575.5050 198.2400 577.5050 ;
        RECT 204.7550 575.5050 206.7550 577.5050 ;
        RECT 204.7550 568.4100 206.7550 570.4100 ;
        RECT 196.2400 568.4100 198.2400 570.4100 ;
        RECT 187.7250 568.4100 189.7250 570.4100 ;
        RECT 179.2100 568.4100 181.2100 570.4100 ;
        RECT 204.7550 561.3150 206.7550 563.3150 ;
        RECT 196.2400 561.3150 198.2400 563.3150 ;
        RECT 187.7250 561.3150 189.7250 563.3150 ;
        RECT 179.2100 561.3150 181.2100 563.3150 ;
        RECT 179.2100 582.6000 181.2100 584.6000 ;
        RECT 187.7250 582.6000 189.7250 584.6000 ;
        RECT 196.2400 582.6000 198.2400 584.6000 ;
        RECT 204.7550 582.6000 206.7550 584.6000 ;
        RECT 179.2100 589.6950 181.2100 591.6950 ;
        RECT 187.7250 589.6950 189.7250 591.6950 ;
        RECT 196.2400 589.6950 198.2400 591.6950 ;
        RECT 204.7550 589.6950 206.7550 591.6950 ;
        RECT 145.1500 610.9800 147.1500 612.9800 ;
        RECT 153.6650 610.9800 155.6650 612.9800 ;
        RECT 162.1800 610.9800 164.1800 612.9800 ;
        RECT 170.6950 610.9800 172.6950 612.9800 ;
        RECT 170.6950 603.8850 172.6950 605.8850 ;
        RECT 162.1800 603.8850 164.1800 605.8850 ;
        RECT 153.6650 603.8850 155.6650 605.8850 ;
        RECT 145.1500 603.8850 147.1500 605.8850 ;
        RECT 170.6950 596.7900 172.6950 598.7900 ;
        RECT 162.1800 596.7900 164.1800 598.7900 ;
        RECT 153.6650 596.7900 155.6650 598.7900 ;
        RECT 145.1500 596.7900 147.1500 598.7900 ;
        RECT 145.1500 618.0750 147.1500 620.0750 ;
        RECT 153.6650 618.0750 155.6650 620.0750 ;
        RECT 162.1800 618.0750 164.1800 620.0750 ;
        RECT 170.6950 618.0750 172.6950 620.0750 ;
        RECT 145.1500 625.1700 147.1500 627.1700 ;
        RECT 153.6650 625.1700 155.6650 627.1700 ;
        RECT 162.1800 625.1700 164.1800 627.1700 ;
        RECT 170.6950 625.1700 172.6950 627.1700 ;
        RECT 179.2100 610.9800 181.2100 612.9800 ;
        RECT 187.7250 610.9800 189.7250 612.9800 ;
        RECT 196.2400 610.9800 198.2400 612.9800 ;
        RECT 204.7550 610.9800 206.7550 612.9800 ;
        RECT 204.7550 603.8850 206.7550 605.8850 ;
        RECT 196.2400 603.8850 198.2400 605.8850 ;
        RECT 187.7250 603.8850 189.7250 605.8850 ;
        RECT 179.2100 603.8850 181.2100 605.8850 ;
        RECT 204.7550 596.7900 206.7550 598.7900 ;
        RECT 196.2400 596.7900 198.2400 598.7900 ;
        RECT 187.7250 596.7900 189.7250 598.7900 ;
        RECT 179.2100 596.7900 181.2100 598.7900 ;
        RECT 179.2100 618.0750 181.2100 620.0750 ;
        RECT 187.7250 618.0750 189.7250 620.0750 ;
        RECT 196.2400 618.0750 198.2400 620.0750 ;
        RECT 204.7550 618.0750 206.7550 620.0750 ;
        RECT 179.2100 625.1700 181.2100 627.1700 ;
        RECT 187.7250 625.1700 189.7250 627.1700 ;
        RECT 196.2400 625.1700 198.2400 627.1700 ;
        RECT 204.7550 625.1700 206.7550 627.1700 ;
        RECT 213.2700 575.5050 215.2700 577.5050 ;
        RECT 221.7850 575.5050 223.7850 577.5050 ;
        RECT 230.3000 575.5050 232.3000 577.5050 ;
        RECT 238.8150 575.5050 240.8150 577.5050 ;
        RECT 238.8150 568.4100 240.8150 570.4100 ;
        RECT 230.3000 568.4100 232.3000 570.4100 ;
        RECT 221.7850 568.4100 223.7850 570.4100 ;
        RECT 213.2700 568.4100 215.2700 570.4100 ;
        RECT 238.8150 561.3150 240.8150 563.3150 ;
        RECT 230.3000 561.3150 232.3000 563.3150 ;
        RECT 221.7850 561.3150 223.7850 563.3150 ;
        RECT 213.2700 561.3150 215.2700 563.3150 ;
        RECT 213.2700 582.6000 215.2700 584.6000 ;
        RECT 221.7850 582.6000 223.7850 584.6000 ;
        RECT 230.3000 582.6000 232.3000 584.6000 ;
        RECT 238.8150 582.6000 240.8150 584.6000 ;
        RECT 213.2700 589.6950 215.2700 591.6950 ;
        RECT 221.7850 589.6950 223.7850 591.6950 ;
        RECT 230.3000 589.6950 232.3000 591.6950 ;
        RECT 238.8150 589.6950 240.8150 591.6950 ;
        RECT 247.3300 575.5050 249.3300 577.5050 ;
        RECT 255.8450 575.5050 257.8450 577.5050 ;
        RECT 264.3600 575.5050 266.3600 577.5050 ;
        RECT 272.8750 575.5050 274.8750 577.5050 ;
        RECT 272.8750 568.4100 274.8750 570.4100 ;
        RECT 264.3600 568.4100 266.3600 570.4100 ;
        RECT 255.8450 568.4100 257.8450 570.4100 ;
        RECT 247.3300 568.4100 249.3300 570.4100 ;
        RECT 272.8750 561.3150 274.8750 563.3150 ;
        RECT 264.3600 561.3150 266.3600 563.3150 ;
        RECT 255.8450 561.3150 257.8450 563.3150 ;
        RECT 247.3300 561.3150 249.3300 563.3150 ;
        RECT 247.3300 582.6000 249.3300 584.6000 ;
        RECT 255.8450 582.6000 257.8450 584.6000 ;
        RECT 264.3600 582.6000 266.3600 584.6000 ;
        RECT 272.8750 582.6000 274.8750 584.6000 ;
        RECT 247.3300 589.6950 249.3300 591.6950 ;
        RECT 255.8450 589.6950 257.8450 591.6950 ;
        RECT 264.3600 589.6950 266.3600 591.6950 ;
        RECT 272.8750 589.6950 274.8750 591.6950 ;
        RECT 213.2700 610.9800 215.2700 612.9800 ;
        RECT 221.7850 610.9800 223.7850 612.9800 ;
        RECT 230.3000 610.9800 232.3000 612.9800 ;
        RECT 238.8150 610.9800 240.8150 612.9800 ;
        RECT 238.8150 603.8850 240.8150 605.8850 ;
        RECT 230.3000 603.8850 232.3000 605.8850 ;
        RECT 221.7850 603.8850 223.7850 605.8850 ;
        RECT 213.2700 603.8850 215.2700 605.8850 ;
        RECT 238.8150 596.7900 240.8150 598.7900 ;
        RECT 230.3000 596.7900 232.3000 598.7900 ;
        RECT 221.7850 596.7900 223.7850 598.7900 ;
        RECT 213.2700 596.7900 215.2700 598.7900 ;
        RECT 213.2700 618.0750 215.2700 620.0750 ;
        RECT 221.7850 618.0750 223.7850 620.0750 ;
        RECT 230.3000 618.0750 232.3000 620.0750 ;
        RECT 238.8150 618.0750 240.8150 620.0750 ;
        RECT 213.2700 625.1700 215.2700 627.1700 ;
        RECT 221.7850 625.1700 223.7850 627.1700 ;
        RECT 230.3000 625.1700 232.3000 627.1700 ;
        RECT 238.8150 625.1700 240.8150 627.1700 ;
        RECT 247.3300 610.9800 249.3300 612.9800 ;
        RECT 255.8450 610.9800 257.8450 612.9800 ;
        RECT 264.3600 610.9800 266.3600 612.9800 ;
        RECT 272.8750 610.9800 274.8750 612.9800 ;
        RECT 272.8750 603.8850 274.8750 605.8850 ;
        RECT 264.3600 603.8850 266.3600 605.8850 ;
        RECT 255.8450 603.8850 257.8450 605.8850 ;
        RECT 247.3300 603.8850 249.3300 605.8850 ;
        RECT 272.8750 596.7900 274.8750 598.7900 ;
        RECT 264.3600 596.7900 266.3600 598.7900 ;
        RECT 255.8450 596.7900 257.8450 598.7900 ;
        RECT 247.3300 596.7900 249.3300 598.7900 ;
        RECT 247.3300 618.0750 249.3300 620.0750 ;
        RECT 255.8450 618.0750 257.8450 620.0750 ;
        RECT 264.3600 618.0750 266.3600 620.0750 ;
        RECT 272.8750 618.0750 274.8750 620.0750 ;
        RECT 247.3300 625.1700 249.3300 627.1700 ;
        RECT 255.8450 625.1700 257.8450 627.1700 ;
        RECT 264.3600 625.1700 266.3600 627.1700 ;
        RECT 272.8750 625.1700 274.8750 627.1700 ;
        RECT 145.1500 646.4550 147.1500 648.4550 ;
        RECT 153.6650 646.4550 155.6650 648.4550 ;
        RECT 162.1800 646.4550 164.1800 648.4550 ;
        RECT 170.6950 646.4550 172.6950 648.4550 ;
        RECT 170.6950 639.3600 172.6950 641.3600 ;
        RECT 162.1800 639.3600 164.1800 641.3600 ;
        RECT 153.6650 639.3600 155.6650 641.3600 ;
        RECT 145.1500 639.3600 147.1500 641.3600 ;
        RECT 170.6950 632.2650 172.6950 634.2650 ;
        RECT 162.1800 632.2650 164.1800 634.2650 ;
        RECT 153.6650 632.2650 155.6650 634.2650 ;
        RECT 145.1500 632.2650 147.1500 634.2650 ;
        RECT 145.1500 653.5500 147.1500 655.5500 ;
        RECT 153.6650 653.5500 155.6650 655.5500 ;
        RECT 162.1800 653.5500 164.1800 655.5500 ;
        RECT 170.6950 653.5500 172.6950 655.5500 ;
        RECT 145.1500 660.6450 147.1500 662.6450 ;
        RECT 153.6650 660.6450 155.6650 662.6450 ;
        RECT 162.1800 660.6450 164.1800 662.6450 ;
        RECT 170.6950 660.6450 172.6950 662.6450 ;
        RECT 179.2100 646.4550 181.2100 648.4550 ;
        RECT 187.7250 646.4550 189.7250 648.4550 ;
        RECT 196.2400 646.4550 198.2400 648.4550 ;
        RECT 204.7550 646.4550 206.7550 648.4550 ;
        RECT 204.7550 639.3600 206.7550 641.3600 ;
        RECT 196.2400 639.3600 198.2400 641.3600 ;
        RECT 187.7250 639.3600 189.7250 641.3600 ;
        RECT 179.2100 639.3600 181.2100 641.3600 ;
        RECT 204.7550 632.2650 206.7550 634.2650 ;
        RECT 196.2400 632.2650 198.2400 634.2650 ;
        RECT 187.7250 632.2650 189.7250 634.2650 ;
        RECT 179.2100 632.2650 181.2100 634.2650 ;
        RECT 179.2100 653.5500 181.2100 655.5500 ;
        RECT 187.7250 653.5500 189.7250 655.5500 ;
        RECT 196.2400 653.5500 198.2400 655.5500 ;
        RECT 204.7550 653.5500 206.7550 655.5500 ;
        RECT 179.2100 660.6450 181.2100 662.6450 ;
        RECT 187.7250 660.6450 189.7250 662.6450 ;
        RECT 196.2400 660.6450 198.2400 662.6450 ;
        RECT 204.7550 660.6450 206.7550 662.6450 ;
        RECT 170.6950 674.8350 172.6950 676.8350 ;
        RECT 162.1800 674.8350 164.1800 676.8350 ;
        RECT 153.6650 674.8350 155.6650 676.8350 ;
        RECT 145.1500 674.8350 147.1500 676.8350 ;
        RECT 170.6950 667.7400 172.6950 669.7400 ;
        RECT 162.1800 667.7400 164.1800 669.7400 ;
        RECT 153.6650 667.7400 155.6650 669.7400 ;
        RECT 145.1500 667.7400 147.1500 669.7400 ;
        RECT 187.7250 674.8350 189.7250 676.8350 ;
        RECT 179.2100 674.8350 181.2100 676.8350 ;
        RECT 204.7550 667.7400 206.7550 669.7400 ;
        RECT 196.2400 667.7400 198.2400 669.7400 ;
        RECT 187.7250 667.7400 189.7250 669.7400 ;
        RECT 179.2100 667.7400 181.2100 669.7400 ;
        RECT 196.2400 674.8350 198.2400 676.8350 ;
        RECT 204.7550 674.8350 206.7550 676.8350 ;
        RECT 213.2700 646.4550 215.2700 648.4550 ;
        RECT 221.7850 646.4550 223.7850 648.4550 ;
        RECT 230.3000 646.4550 232.3000 648.4550 ;
        RECT 238.8150 646.4550 240.8150 648.4550 ;
        RECT 238.8150 639.3600 240.8150 641.3600 ;
        RECT 230.3000 639.3600 232.3000 641.3600 ;
        RECT 221.7850 639.3600 223.7850 641.3600 ;
        RECT 213.2700 639.3600 215.2700 641.3600 ;
        RECT 238.8150 632.2650 240.8150 634.2650 ;
        RECT 230.3000 632.2650 232.3000 634.2650 ;
        RECT 221.7850 632.2650 223.7850 634.2650 ;
        RECT 213.2700 632.2650 215.2700 634.2650 ;
        RECT 213.2700 653.5500 215.2700 655.5500 ;
        RECT 221.7850 653.5500 223.7850 655.5500 ;
        RECT 230.3000 653.5500 232.3000 655.5500 ;
        RECT 238.8150 653.5500 240.8150 655.5500 ;
        RECT 213.2700 660.6450 215.2700 662.6450 ;
        RECT 221.7850 660.6450 223.7850 662.6450 ;
        RECT 230.3000 660.6450 232.3000 662.6450 ;
        RECT 238.8150 660.6450 240.8150 662.6450 ;
        RECT 247.3300 646.4550 249.3300 648.4550 ;
        RECT 255.8450 646.4550 257.8450 648.4550 ;
        RECT 264.3600 646.4550 266.3600 648.4550 ;
        RECT 272.8750 646.4550 274.8750 648.4550 ;
        RECT 272.8750 639.3600 274.8750 641.3600 ;
        RECT 264.3600 639.3600 266.3600 641.3600 ;
        RECT 255.8450 639.3600 257.8450 641.3600 ;
        RECT 247.3300 639.3600 249.3300 641.3600 ;
        RECT 272.8750 632.2650 274.8750 634.2650 ;
        RECT 264.3600 632.2650 266.3600 634.2650 ;
        RECT 255.8450 632.2650 257.8450 634.2650 ;
        RECT 247.3300 632.2650 249.3300 634.2650 ;
        RECT 247.3300 653.5500 249.3300 655.5500 ;
        RECT 255.8450 653.5500 257.8450 655.5500 ;
        RECT 264.3600 653.5500 266.3600 655.5500 ;
        RECT 272.8750 653.5500 274.8750 655.5500 ;
        RECT 247.3300 660.6450 249.3300 662.6450 ;
        RECT 255.8450 660.6450 257.8450 662.6450 ;
        RECT 264.3600 660.6450 266.3600 662.6450 ;
        RECT 272.8750 660.6450 274.8750 662.6450 ;
        RECT 238.8150 674.8350 240.8150 676.8350 ;
        RECT 230.3000 674.8350 232.3000 676.8350 ;
        RECT 221.7850 674.8350 223.7850 676.8350 ;
        RECT 213.2700 674.8350 215.2700 676.8350 ;
        RECT 238.8150 667.7400 240.8150 669.7400 ;
        RECT 230.3000 667.7400 232.3000 669.7400 ;
        RECT 221.7850 667.7400 223.7850 669.7400 ;
        RECT 213.2700 667.7400 215.2700 669.7400 ;
        RECT 255.8450 674.8350 257.8450 676.8350 ;
        RECT 247.3300 674.8350 249.3300 676.8350 ;
        RECT 272.8750 667.7400 274.8750 669.7400 ;
        RECT 264.3600 667.7400 266.3600 669.7400 ;
        RECT 255.8450 667.7400 257.8450 669.7400 ;
        RECT 247.3300 667.7400 249.3300 669.7400 ;
        RECT 264.3600 674.8350 266.3600 676.8350 ;
        RECT 272.8750 674.8350 274.8750 676.8350 ;
        RECT 6.0000 717.4050 8.0000 719.4050 ;
        RECT 6.0000 710.3100 8.0000 712.3100 ;
        RECT 6.0000 703.2150 8.0000 705.2150 ;
        RECT 6.0000 731.5950 8.0000 733.5950 ;
        RECT 6.0000 724.5000 8.0000 726.5000 ;
        RECT 6.0000 738.6900 8.0000 740.6900 ;
        RECT 6.0000 745.7850 8.0000 747.7850 ;
        RECT 6.0000 759.9750 8.0000 761.9750 ;
        RECT 6.0000 752.8800 8.0000 754.8800 ;
        RECT 6.0000 767.0700 8.0000 769.0700 ;
        RECT 6.0000 781.2600 8.0000 783.2600 ;
        RECT 6.0000 774.1650 8.0000 776.1650 ;
        RECT 6.0000 795.4500 8.0000 797.4500 ;
        RECT 6.0000 788.3550 8.0000 790.3550 ;
        RECT 6.0000 802.5450 8.0000 804.5450 ;
        RECT 6.0000 809.6400 8.0000 811.6400 ;
        RECT 6.0000 816.7350 8.0000 818.7350 ;
        RECT 6.0000 830.9250 8.0000 832.9250 ;
        RECT 6.0000 823.8300 8.0000 825.8300 ;
        RECT 281.3900 575.5050 283.3900 577.5050 ;
        RECT 289.9050 575.5050 291.9050 577.5050 ;
        RECT 298.4200 575.5050 300.4200 577.5050 ;
        RECT 306.9350 575.5050 308.9350 577.5050 ;
        RECT 306.9350 568.4100 308.9350 570.4100 ;
        RECT 298.4200 568.4100 300.4200 570.4100 ;
        RECT 289.9050 568.4100 291.9050 570.4100 ;
        RECT 281.3900 568.4100 283.3900 570.4100 ;
        RECT 306.9350 561.3150 308.9350 563.3150 ;
        RECT 298.4200 561.3150 300.4200 563.3150 ;
        RECT 289.9050 561.3150 291.9050 563.3150 ;
        RECT 281.3900 561.3150 283.3900 563.3150 ;
        RECT 281.3900 582.6000 283.3900 584.6000 ;
        RECT 289.9050 582.6000 291.9050 584.6000 ;
        RECT 298.4200 582.6000 300.4200 584.6000 ;
        RECT 306.9350 582.6000 308.9350 584.6000 ;
        RECT 281.3900 589.6950 283.3900 591.6950 ;
        RECT 289.9050 589.6950 291.9050 591.6950 ;
        RECT 298.4200 589.6950 300.4200 591.6950 ;
        RECT 306.9350 589.6950 308.9350 591.6950 ;
        RECT 344.0000 575.5050 346.0000 577.5050 ;
        RECT 315.4500 575.5050 317.4500 577.5050 ;
        RECT 323.9650 575.5050 325.9650 577.5050 ;
        RECT 323.9650 568.4100 325.9650 570.4100 ;
        RECT 315.4500 568.4100 317.4500 570.4100 ;
        RECT 323.9650 561.3150 325.9650 563.3150 ;
        RECT 315.4500 561.3150 317.4500 563.3150 ;
        RECT 344.0000 568.4100 346.0000 570.4100 ;
        RECT 344.0000 561.3150 346.0000 563.3150 ;
        RECT 323.9650 589.6950 325.9650 591.6950 ;
        RECT 315.4500 589.6950 317.4500 591.6950 ;
        RECT 323.9650 582.6000 325.9650 584.6000 ;
        RECT 315.4500 582.6000 317.4500 584.6000 ;
        RECT 344.0000 589.6950 346.0000 591.6950 ;
        RECT 344.0000 582.6000 346.0000 584.6000 ;
        RECT 281.3900 610.9800 283.3900 612.9800 ;
        RECT 289.9050 610.9800 291.9050 612.9800 ;
        RECT 298.4200 610.9800 300.4200 612.9800 ;
        RECT 306.9350 610.9800 308.9350 612.9800 ;
        RECT 306.9350 603.8850 308.9350 605.8850 ;
        RECT 298.4200 603.8850 300.4200 605.8850 ;
        RECT 289.9050 603.8850 291.9050 605.8850 ;
        RECT 281.3900 603.8850 283.3900 605.8850 ;
        RECT 306.9350 596.7900 308.9350 598.7900 ;
        RECT 298.4200 596.7900 300.4200 598.7900 ;
        RECT 289.9050 596.7900 291.9050 598.7900 ;
        RECT 281.3900 596.7900 283.3900 598.7900 ;
        RECT 281.3900 618.0750 283.3900 620.0750 ;
        RECT 289.9050 618.0750 291.9050 620.0750 ;
        RECT 298.4200 618.0750 300.4200 620.0750 ;
        RECT 306.9350 618.0750 308.9350 620.0750 ;
        RECT 281.3900 625.1700 283.3900 627.1700 ;
        RECT 289.9050 625.1700 291.9050 627.1700 ;
        RECT 298.4200 625.1700 300.4200 627.1700 ;
        RECT 306.9350 625.1700 308.9350 627.1700 ;
        RECT 344.0000 610.9800 346.0000 612.9800 ;
        RECT 315.4500 610.9800 317.4500 612.9800 ;
        RECT 323.9650 610.9800 325.9650 612.9800 ;
        RECT 323.9650 603.8850 325.9650 605.8850 ;
        RECT 315.4500 603.8850 317.4500 605.8850 ;
        RECT 323.9650 596.7900 325.9650 598.7900 ;
        RECT 315.4500 596.7900 317.4500 598.7900 ;
        RECT 344.0000 603.8850 346.0000 605.8850 ;
        RECT 344.0000 596.7900 346.0000 598.7900 ;
        RECT 323.9650 618.0750 325.9650 620.0750 ;
        RECT 315.4500 618.0750 317.4500 620.0750 ;
        RECT 315.4500 625.1700 317.4500 627.1700 ;
        RECT 323.9650 625.1700 325.9650 627.1700 ;
        RECT 344.0000 625.1700 346.0000 627.1700 ;
        RECT 344.0000 618.0750 346.0000 620.0750 ;
        RECT 394.0000 575.5050 396.0000 577.5050 ;
        RECT 414.1500 575.5050 416.1500 577.5050 ;
        RECT 394.0000 568.4100 396.0000 570.4100 ;
        RECT 394.0000 561.3150 396.0000 563.3150 ;
        RECT 414.1500 568.4100 416.1500 570.4100 ;
        RECT 414.1500 561.3150 416.1500 563.3150 ;
        RECT 394.0000 582.6000 396.0000 584.6000 ;
        RECT 394.0000 589.6950 396.0000 591.6950 ;
        RECT 414.1500 582.6000 416.1500 584.6000 ;
        RECT 414.1500 589.6950 416.1500 591.6950 ;
        RECT 394.0000 610.9800 396.0000 612.9800 ;
        RECT 414.1500 610.9800 416.1500 612.9800 ;
        RECT 394.0000 596.7900 396.0000 598.7900 ;
        RECT 394.0000 603.8850 396.0000 605.8850 ;
        RECT 414.1500 596.7900 416.1500 598.7900 ;
        RECT 414.1500 603.8850 416.1500 605.8850 ;
        RECT 394.0000 625.1700 396.0000 627.1700 ;
        RECT 394.0000 618.0750 396.0000 620.0750 ;
        RECT 414.1500 625.1700 416.1500 627.1700 ;
        RECT 414.1500 618.0750 416.1500 620.0750 ;
        RECT 281.3900 646.4550 283.3900 648.4550 ;
        RECT 289.9050 646.4550 291.9050 648.4550 ;
        RECT 298.4200 646.4550 300.4200 648.4550 ;
        RECT 306.9350 646.4550 308.9350 648.4550 ;
        RECT 306.9350 639.3600 308.9350 641.3600 ;
        RECT 298.4200 639.3600 300.4200 641.3600 ;
        RECT 289.9050 639.3600 291.9050 641.3600 ;
        RECT 281.3900 639.3600 283.3900 641.3600 ;
        RECT 306.9350 632.2650 308.9350 634.2650 ;
        RECT 298.4200 632.2650 300.4200 634.2650 ;
        RECT 289.9050 632.2650 291.9050 634.2650 ;
        RECT 281.3900 632.2650 283.3900 634.2650 ;
        RECT 281.3900 653.5500 283.3900 655.5500 ;
        RECT 289.9050 653.5500 291.9050 655.5500 ;
        RECT 298.4200 653.5500 300.4200 655.5500 ;
        RECT 306.9350 653.5500 308.9350 655.5500 ;
        RECT 281.3900 660.6450 283.3900 662.6450 ;
        RECT 289.9050 660.6450 291.9050 662.6450 ;
        RECT 298.4200 660.6450 300.4200 662.6450 ;
        RECT 306.9350 660.6450 308.9350 662.6450 ;
        RECT 344.0000 646.4550 346.0000 648.4550 ;
        RECT 315.4500 646.4550 317.4500 648.4550 ;
        RECT 323.9650 646.4550 325.9650 648.4550 ;
        RECT 315.4500 639.3600 317.4500 641.3600 ;
        RECT 323.9650 632.2650 325.9650 634.2650 ;
        RECT 315.4500 632.2650 317.4500 634.2650 ;
        RECT 323.9650 639.3600 325.9650 641.3600 ;
        RECT 344.0000 632.2650 346.0000 634.2650 ;
        RECT 344.0000 639.3600 346.0000 641.3600 ;
        RECT 323.9650 660.6450 325.9650 662.6450 ;
        RECT 315.4500 660.6450 317.4500 662.6450 ;
        RECT 323.9650 653.5500 325.9650 655.5500 ;
        RECT 315.4500 653.5500 317.4500 655.5500 ;
        RECT 344.0000 653.5500 346.0000 655.5500 ;
        RECT 344.0000 660.6450 346.0000 662.6450 ;
        RECT 281.3900 667.7400 283.3900 669.7400 ;
        RECT 289.9050 667.7400 291.9050 669.7400 ;
        RECT 298.4200 667.7400 300.4200 669.7400 ;
        RECT 306.9350 667.7400 308.9350 669.7400 ;
        RECT 281.3900 674.8350 283.3900 676.8350 ;
        RECT 289.9050 674.8350 291.9050 676.8350 ;
        RECT 298.4200 674.8350 300.4200 676.8350 ;
        RECT 306.9350 674.8350 308.9350 676.8350 ;
        RECT 344.0000 681.9300 346.0000 683.9300 ;
        RECT 323.9650 667.7400 325.9650 669.7400 ;
        RECT 315.4500 667.7400 317.4500 669.7400 ;
        RECT 315.4500 674.8350 317.4500 676.8350 ;
        RECT 323.9650 674.8350 325.9650 676.8350 ;
        RECT 344.0000 667.7400 346.0000 669.7400 ;
        RECT 344.0000 674.8350 346.0000 676.8350 ;
        RECT 344.0000 689.0250 346.0000 691.0250 ;
        RECT 394.0000 646.4550 396.0000 648.4550 ;
        RECT 414.1500 646.4550 416.1500 648.4550 ;
        RECT 394.0000 639.3600 396.0000 641.3600 ;
        RECT 394.0000 632.2650 396.0000 634.2650 ;
        RECT 414.1500 639.3600 416.1500 641.3600 ;
        RECT 414.1500 632.2650 416.1500 634.2650 ;
        RECT 394.0000 653.5500 396.0000 655.5500 ;
        RECT 394.0000 660.6450 396.0000 662.6450 ;
        RECT 414.1500 653.5500 416.1500 655.5500 ;
        RECT 414.1500 660.6450 416.1500 662.6450 ;
        RECT 394.0000 681.9300 396.0000 683.9300 ;
        RECT 414.1500 681.9300 416.1500 683.9300 ;
        RECT 394.0000 674.8350 396.0000 676.8350 ;
        RECT 394.0000 667.7400 396.0000 669.7400 ;
        RECT 414.1500 674.8350 416.1500 676.8350 ;
        RECT 414.1500 667.7400 416.1500 669.7400 ;
        RECT 394.0000 696.1200 396.0000 698.1200 ;
        RECT 394.0000 689.0250 396.0000 691.0250 ;
        RECT 414.1500 696.1200 416.1500 698.1200 ;
        RECT 414.1500 689.0250 416.1500 691.0250 ;
        RECT 454.9000 561.3150 456.9000 563.3150 ;
        RECT 454.9000 568.4100 456.9000 570.4100 ;
        RECT 454.9000 575.5050 456.9000 577.5050 ;
        RECT 454.9000 582.6000 456.9000 584.6000 ;
        RECT 454.9000 589.6950 456.9000 591.6950 ;
        RECT 422.3000 575.5050 424.3000 577.5050 ;
        RECT 430.4500 575.5050 432.4500 577.5050 ;
        RECT 438.6000 575.5050 440.6000 577.5050 ;
        RECT 446.7500 575.5050 448.7500 577.5050 ;
        RECT 446.7500 568.4100 448.7500 570.4100 ;
        RECT 438.6000 568.4100 440.6000 570.4100 ;
        RECT 430.4500 568.4100 432.4500 570.4100 ;
        RECT 422.3000 568.4100 424.3000 570.4100 ;
        RECT 446.7500 561.3150 448.7500 563.3150 ;
        RECT 438.6000 561.3150 440.6000 563.3150 ;
        RECT 430.4500 561.3150 432.4500 563.3150 ;
        RECT 422.3000 561.3150 424.3000 563.3150 ;
        RECT 422.3000 582.6000 424.3000 584.6000 ;
        RECT 430.4500 582.6000 432.4500 584.6000 ;
        RECT 438.6000 582.6000 440.6000 584.6000 ;
        RECT 446.7500 582.6000 448.7500 584.6000 ;
        RECT 422.3000 589.6950 424.3000 591.6950 ;
        RECT 430.4500 589.6950 432.4500 591.6950 ;
        RECT 438.6000 589.6950 440.6000 591.6950 ;
        RECT 446.7500 589.6950 448.7500 591.6950 ;
        RECT 463.0500 575.5050 465.0500 577.5050 ;
        RECT 471.2000 575.5050 473.2000 577.5050 ;
        RECT 479.3500 575.5050 481.3500 577.5050 ;
        RECT 487.5000 575.5050 489.5000 577.5050 ;
        RECT 487.5000 568.4100 489.5000 570.4100 ;
        RECT 479.3500 568.4100 481.3500 570.4100 ;
        RECT 471.2000 568.4100 473.2000 570.4100 ;
        RECT 463.0500 568.4100 465.0500 570.4100 ;
        RECT 487.5000 561.3150 489.5000 563.3150 ;
        RECT 479.3500 561.3150 481.3500 563.3150 ;
        RECT 471.2000 561.3150 473.2000 563.3150 ;
        RECT 463.0500 561.3150 465.0500 563.3150 ;
        RECT 463.0500 582.6000 465.0500 584.6000 ;
        RECT 471.2000 582.6000 473.2000 584.6000 ;
        RECT 479.3500 582.6000 481.3500 584.6000 ;
        RECT 487.5000 582.6000 489.5000 584.6000 ;
        RECT 463.0500 589.6950 465.0500 591.6950 ;
        RECT 471.2000 589.6950 473.2000 591.6950 ;
        RECT 479.3500 589.6950 481.3500 591.6950 ;
        RECT 487.5000 589.6950 489.5000 591.6950 ;
        RECT 454.9000 596.7900 456.9000 598.7900 ;
        RECT 454.9000 603.8850 456.9000 605.8850 ;
        RECT 454.9000 610.9800 456.9000 612.9800 ;
        RECT 454.9000 618.0750 456.9000 620.0750 ;
        RECT 454.9000 625.1700 456.9000 627.1700 ;
        RECT 422.3000 610.9800 424.3000 612.9800 ;
        RECT 430.4500 610.9800 432.4500 612.9800 ;
        RECT 438.6000 610.9800 440.6000 612.9800 ;
        RECT 446.7500 610.9800 448.7500 612.9800 ;
        RECT 446.7500 603.8850 448.7500 605.8850 ;
        RECT 438.6000 603.8850 440.6000 605.8850 ;
        RECT 430.4500 603.8850 432.4500 605.8850 ;
        RECT 422.3000 603.8850 424.3000 605.8850 ;
        RECT 446.7500 596.7900 448.7500 598.7900 ;
        RECT 438.6000 596.7900 440.6000 598.7900 ;
        RECT 430.4500 596.7900 432.4500 598.7900 ;
        RECT 422.3000 596.7900 424.3000 598.7900 ;
        RECT 422.3000 618.0750 424.3000 620.0750 ;
        RECT 430.4500 618.0750 432.4500 620.0750 ;
        RECT 438.6000 618.0750 440.6000 620.0750 ;
        RECT 446.7500 618.0750 448.7500 620.0750 ;
        RECT 422.3000 625.1700 424.3000 627.1700 ;
        RECT 430.4500 625.1700 432.4500 627.1700 ;
        RECT 438.6000 625.1700 440.6000 627.1700 ;
        RECT 446.7500 625.1700 448.7500 627.1700 ;
        RECT 463.0500 610.9800 465.0500 612.9800 ;
        RECT 471.2000 610.9800 473.2000 612.9800 ;
        RECT 479.3500 610.9800 481.3500 612.9800 ;
        RECT 487.5000 610.9800 489.5000 612.9800 ;
        RECT 487.5000 603.8850 489.5000 605.8850 ;
        RECT 479.3500 603.8850 481.3500 605.8850 ;
        RECT 471.2000 603.8850 473.2000 605.8850 ;
        RECT 463.0500 603.8850 465.0500 605.8850 ;
        RECT 487.5000 596.7900 489.5000 598.7900 ;
        RECT 479.3500 596.7900 481.3500 598.7900 ;
        RECT 471.2000 596.7900 473.2000 598.7900 ;
        RECT 463.0500 596.7900 465.0500 598.7900 ;
        RECT 463.0500 618.0750 465.0500 620.0750 ;
        RECT 471.2000 618.0750 473.2000 620.0750 ;
        RECT 479.3500 618.0750 481.3500 620.0750 ;
        RECT 487.5000 618.0750 489.5000 620.0750 ;
        RECT 463.0500 625.1700 465.0500 627.1700 ;
        RECT 471.2000 625.1700 473.2000 627.1700 ;
        RECT 479.3500 625.1700 481.3500 627.1700 ;
        RECT 487.5000 625.1700 489.5000 627.1700 ;
        RECT 495.6500 575.5050 497.6500 577.5050 ;
        RECT 503.8000 575.5050 505.8000 577.5050 ;
        RECT 511.9500 575.5050 513.9500 577.5050 ;
        RECT 520.1000 575.5050 522.1000 577.5050 ;
        RECT 520.1000 568.4100 522.1000 570.4100 ;
        RECT 511.9500 568.4100 513.9500 570.4100 ;
        RECT 503.8000 568.4100 505.8000 570.4100 ;
        RECT 495.6500 568.4100 497.6500 570.4100 ;
        RECT 520.1000 561.3150 522.1000 563.3150 ;
        RECT 511.9500 561.3150 513.9500 563.3150 ;
        RECT 503.8000 561.3150 505.8000 563.3150 ;
        RECT 495.6500 561.3150 497.6500 563.3150 ;
        RECT 495.6500 582.6000 497.6500 584.6000 ;
        RECT 503.8000 582.6000 505.8000 584.6000 ;
        RECT 511.9500 582.6000 513.9500 584.6000 ;
        RECT 520.1000 582.6000 522.1000 584.6000 ;
        RECT 495.6500 589.6950 497.6500 591.6950 ;
        RECT 503.8000 589.6950 505.8000 591.6950 ;
        RECT 511.9500 589.6950 513.9500 591.6950 ;
        RECT 520.1000 589.6950 522.1000 591.6950 ;
        RECT 528.2500 575.5050 530.2500 577.5050 ;
        RECT 536.4000 575.5050 538.4000 577.5050 ;
        RECT 544.5500 575.5050 546.5500 577.5050 ;
        RECT 552.7000 575.5050 554.7000 577.5050 ;
        RECT 552.7000 568.4100 554.7000 570.4100 ;
        RECT 544.5500 568.4100 546.5500 570.4100 ;
        RECT 536.4000 568.4100 538.4000 570.4100 ;
        RECT 528.2500 568.4100 530.2500 570.4100 ;
        RECT 552.7000 561.3150 554.7000 563.3150 ;
        RECT 544.5500 561.3150 546.5500 563.3150 ;
        RECT 536.4000 561.3150 538.4000 563.3150 ;
        RECT 528.2500 561.3150 530.2500 563.3150 ;
        RECT 528.2500 582.6000 530.2500 584.6000 ;
        RECT 536.4000 582.6000 538.4000 584.6000 ;
        RECT 544.5500 582.6000 546.5500 584.6000 ;
        RECT 552.7000 582.6000 554.7000 584.6000 ;
        RECT 528.2500 589.6950 530.2500 591.6950 ;
        RECT 536.4000 589.6950 538.4000 591.6950 ;
        RECT 544.5500 589.6950 546.5500 591.6950 ;
        RECT 552.7000 589.6950 554.7000 591.6950 ;
        RECT 495.6500 610.9800 497.6500 612.9800 ;
        RECT 503.8000 610.9800 505.8000 612.9800 ;
        RECT 511.9500 610.9800 513.9500 612.9800 ;
        RECT 520.1000 610.9800 522.1000 612.9800 ;
        RECT 520.1000 603.8850 522.1000 605.8850 ;
        RECT 511.9500 603.8850 513.9500 605.8850 ;
        RECT 503.8000 603.8850 505.8000 605.8850 ;
        RECT 495.6500 603.8850 497.6500 605.8850 ;
        RECT 520.1000 596.7900 522.1000 598.7900 ;
        RECT 511.9500 596.7900 513.9500 598.7900 ;
        RECT 503.8000 596.7900 505.8000 598.7900 ;
        RECT 495.6500 596.7900 497.6500 598.7900 ;
        RECT 495.6500 618.0750 497.6500 620.0750 ;
        RECT 503.8000 618.0750 505.8000 620.0750 ;
        RECT 511.9500 618.0750 513.9500 620.0750 ;
        RECT 520.1000 618.0750 522.1000 620.0750 ;
        RECT 495.6500 625.1700 497.6500 627.1700 ;
        RECT 503.8000 625.1700 505.8000 627.1700 ;
        RECT 511.9500 625.1700 513.9500 627.1700 ;
        RECT 520.1000 625.1700 522.1000 627.1700 ;
        RECT 528.2500 610.9800 530.2500 612.9800 ;
        RECT 536.4000 610.9800 538.4000 612.9800 ;
        RECT 544.5500 610.9800 546.5500 612.9800 ;
        RECT 552.7000 610.9800 554.7000 612.9800 ;
        RECT 552.7000 603.8850 554.7000 605.8850 ;
        RECT 544.5500 603.8850 546.5500 605.8850 ;
        RECT 536.4000 603.8850 538.4000 605.8850 ;
        RECT 528.2500 603.8850 530.2500 605.8850 ;
        RECT 552.7000 596.7900 554.7000 598.7900 ;
        RECT 544.5500 596.7900 546.5500 598.7900 ;
        RECT 536.4000 596.7900 538.4000 598.7900 ;
        RECT 528.2500 596.7900 530.2500 598.7900 ;
        RECT 528.2500 618.0750 530.2500 620.0750 ;
        RECT 536.4000 618.0750 538.4000 620.0750 ;
        RECT 544.5500 618.0750 546.5500 620.0750 ;
        RECT 552.7000 618.0750 554.7000 620.0750 ;
        RECT 528.2500 625.1700 530.2500 627.1700 ;
        RECT 536.4000 625.1700 538.4000 627.1700 ;
        RECT 544.5500 625.1700 546.5500 627.1700 ;
        RECT 552.7000 625.1700 554.7000 627.1700 ;
        RECT 454.9000 632.2650 456.9000 634.2650 ;
        RECT 454.9000 639.3600 456.9000 641.3600 ;
        RECT 454.9000 646.4550 456.9000 648.4550 ;
        RECT 454.9000 653.5500 456.9000 655.5500 ;
        RECT 454.9000 660.6450 456.9000 662.6450 ;
        RECT 422.3000 646.4550 424.3000 648.4550 ;
        RECT 430.4500 646.4550 432.4500 648.4550 ;
        RECT 438.6000 646.4550 440.6000 648.4550 ;
        RECT 446.7500 646.4550 448.7500 648.4550 ;
        RECT 446.7500 639.3600 448.7500 641.3600 ;
        RECT 438.6000 639.3600 440.6000 641.3600 ;
        RECT 430.4500 639.3600 432.4500 641.3600 ;
        RECT 422.3000 639.3600 424.3000 641.3600 ;
        RECT 446.7500 632.2650 448.7500 634.2650 ;
        RECT 438.6000 632.2650 440.6000 634.2650 ;
        RECT 430.4500 632.2650 432.4500 634.2650 ;
        RECT 422.3000 632.2650 424.3000 634.2650 ;
        RECT 422.3000 653.5500 424.3000 655.5500 ;
        RECT 430.4500 653.5500 432.4500 655.5500 ;
        RECT 438.6000 653.5500 440.6000 655.5500 ;
        RECT 446.7500 653.5500 448.7500 655.5500 ;
        RECT 422.3000 660.6450 424.3000 662.6450 ;
        RECT 430.4500 660.6450 432.4500 662.6450 ;
        RECT 438.6000 660.6450 440.6000 662.6450 ;
        RECT 446.7500 660.6450 448.7500 662.6450 ;
        RECT 463.0500 646.4550 465.0500 648.4550 ;
        RECT 471.2000 646.4550 473.2000 648.4550 ;
        RECT 479.3500 646.4550 481.3500 648.4550 ;
        RECT 487.5000 646.4550 489.5000 648.4550 ;
        RECT 487.5000 639.3600 489.5000 641.3600 ;
        RECT 479.3500 639.3600 481.3500 641.3600 ;
        RECT 471.2000 639.3600 473.2000 641.3600 ;
        RECT 463.0500 639.3600 465.0500 641.3600 ;
        RECT 487.5000 632.2650 489.5000 634.2650 ;
        RECT 479.3500 632.2650 481.3500 634.2650 ;
        RECT 471.2000 632.2650 473.2000 634.2650 ;
        RECT 463.0500 632.2650 465.0500 634.2650 ;
        RECT 463.0500 653.5500 465.0500 655.5500 ;
        RECT 471.2000 653.5500 473.2000 655.5500 ;
        RECT 479.3500 653.5500 481.3500 655.5500 ;
        RECT 487.5000 653.5500 489.5000 655.5500 ;
        RECT 463.0500 660.6450 465.0500 662.6450 ;
        RECT 471.2000 660.6450 473.2000 662.6450 ;
        RECT 479.3500 660.6450 481.3500 662.6450 ;
        RECT 487.5000 660.6450 489.5000 662.6450 ;
        RECT 454.9000 667.7400 456.9000 669.7400 ;
        RECT 454.9000 674.8350 456.9000 676.8350 ;
        RECT 454.9000 681.9300 456.9000 683.9300 ;
        RECT 454.9000 689.0250 456.9000 691.0250 ;
        RECT 454.9000 696.1200 456.9000 698.1200 ;
        RECT 422.3000 681.9300 424.3000 683.9300 ;
        RECT 430.4500 681.9300 432.4500 683.9300 ;
        RECT 438.6000 681.9300 440.6000 683.9300 ;
        RECT 446.7500 681.9300 448.7500 683.9300 ;
        RECT 446.7500 674.8350 448.7500 676.8350 ;
        RECT 438.6000 674.8350 440.6000 676.8350 ;
        RECT 430.4500 674.8350 432.4500 676.8350 ;
        RECT 422.3000 674.8350 424.3000 676.8350 ;
        RECT 446.7500 667.7400 448.7500 669.7400 ;
        RECT 438.6000 667.7400 440.6000 669.7400 ;
        RECT 430.4500 667.7400 432.4500 669.7400 ;
        RECT 422.3000 667.7400 424.3000 669.7400 ;
        RECT 422.3000 689.0250 424.3000 691.0250 ;
        RECT 430.4500 689.0250 432.4500 691.0250 ;
        RECT 438.6000 689.0250 440.6000 691.0250 ;
        RECT 446.7500 689.0250 448.7500 691.0250 ;
        RECT 422.3000 696.1200 424.3000 698.1200 ;
        RECT 430.4500 696.1200 432.4500 698.1200 ;
        RECT 438.6000 696.1200 440.6000 698.1200 ;
        RECT 446.7500 696.1200 448.7500 698.1200 ;
        RECT 463.0500 681.9300 465.0500 683.9300 ;
        RECT 471.2000 681.9300 473.2000 683.9300 ;
        RECT 479.3500 681.9300 481.3500 683.9300 ;
        RECT 487.5000 681.9300 489.5000 683.9300 ;
        RECT 487.5000 674.8350 489.5000 676.8350 ;
        RECT 479.3500 674.8350 481.3500 676.8350 ;
        RECT 471.2000 674.8350 473.2000 676.8350 ;
        RECT 463.0500 674.8350 465.0500 676.8350 ;
        RECT 487.5000 667.7400 489.5000 669.7400 ;
        RECT 479.3500 667.7400 481.3500 669.7400 ;
        RECT 471.2000 667.7400 473.2000 669.7400 ;
        RECT 463.0500 667.7400 465.0500 669.7400 ;
        RECT 463.0500 689.0250 465.0500 691.0250 ;
        RECT 471.2000 689.0250 473.2000 691.0250 ;
        RECT 479.3500 689.0250 481.3500 691.0250 ;
        RECT 487.5000 689.0250 489.5000 691.0250 ;
        RECT 463.0500 696.1200 465.0500 698.1200 ;
        RECT 471.2000 696.1200 473.2000 698.1200 ;
        RECT 479.3500 696.1200 481.3500 698.1200 ;
        RECT 487.5000 696.1200 489.5000 698.1200 ;
        RECT 495.6500 646.4550 497.6500 648.4550 ;
        RECT 503.8000 646.4550 505.8000 648.4550 ;
        RECT 511.9500 646.4550 513.9500 648.4550 ;
        RECT 520.1000 646.4550 522.1000 648.4550 ;
        RECT 520.1000 639.3600 522.1000 641.3600 ;
        RECT 511.9500 639.3600 513.9500 641.3600 ;
        RECT 503.8000 639.3600 505.8000 641.3600 ;
        RECT 495.6500 639.3600 497.6500 641.3600 ;
        RECT 520.1000 632.2650 522.1000 634.2650 ;
        RECT 511.9500 632.2650 513.9500 634.2650 ;
        RECT 503.8000 632.2650 505.8000 634.2650 ;
        RECT 495.6500 632.2650 497.6500 634.2650 ;
        RECT 495.6500 653.5500 497.6500 655.5500 ;
        RECT 503.8000 653.5500 505.8000 655.5500 ;
        RECT 511.9500 653.5500 513.9500 655.5500 ;
        RECT 520.1000 653.5500 522.1000 655.5500 ;
        RECT 495.6500 660.6450 497.6500 662.6450 ;
        RECT 503.8000 660.6450 505.8000 662.6450 ;
        RECT 511.9500 660.6450 513.9500 662.6450 ;
        RECT 520.1000 660.6450 522.1000 662.6450 ;
        RECT 528.2500 646.4550 530.2500 648.4550 ;
        RECT 536.4000 646.4550 538.4000 648.4550 ;
        RECT 544.5500 646.4550 546.5500 648.4550 ;
        RECT 552.7000 646.4550 554.7000 648.4550 ;
        RECT 552.7000 639.3600 554.7000 641.3600 ;
        RECT 544.5500 639.3600 546.5500 641.3600 ;
        RECT 536.4000 639.3600 538.4000 641.3600 ;
        RECT 528.2500 639.3600 530.2500 641.3600 ;
        RECT 552.7000 632.2650 554.7000 634.2650 ;
        RECT 544.5500 632.2650 546.5500 634.2650 ;
        RECT 536.4000 632.2650 538.4000 634.2650 ;
        RECT 528.2500 632.2650 530.2500 634.2650 ;
        RECT 528.2500 653.5500 530.2500 655.5500 ;
        RECT 536.4000 653.5500 538.4000 655.5500 ;
        RECT 544.5500 653.5500 546.5500 655.5500 ;
        RECT 552.7000 653.5500 554.7000 655.5500 ;
        RECT 528.2500 660.6450 530.2500 662.6450 ;
        RECT 536.4000 660.6450 538.4000 662.6450 ;
        RECT 544.5500 660.6450 546.5500 662.6450 ;
        RECT 552.7000 660.6450 554.7000 662.6450 ;
        RECT 495.6500 681.9300 497.6500 683.9300 ;
        RECT 503.8000 681.9300 505.8000 683.9300 ;
        RECT 511.9500 681.9300 513.9500 683.9300 ;
        RECT 520.1000 681.9300 522.1000 683.9300 ;
        RECT 520.1000 674.8350 522.1000 676.8350 ;
        RECT 511.9500 674.8350 513.9500 676.8350 ;
        RECT 503.8000 674.8350 505.8000 676.8350 ;
        RECT 495.6500 674.8350 497.6500 676.8350 ;
        RECT 520.1000 667.7400 522.1000 669.7400 ;
        RECT 511.9500 667.7400 513.9500 669.7400 ;
        RECT 503.8000 667.7400 505.8000 669.7400 ;
        RECT 495.6500 667.7400 497.6500 669.7400 ;
        RECT 495.6500 689.0250 497.6500 691.0250 ;
        RECT 503.8000 689.0250 505.8000 691.0250 ;
        RECT 511.9500 689.0250 513.9500 691.0250 ;
        RECT 520.1000 689.0250 522.1000 691.0250 ;
        RECT 495.6500 696.1200 497.6500 698.1200 ;
        RECT 503.8000 696.1200 505.8000 698.1200 ;
        RECT 511.9500 696.1200 513.9500 698.1200 ;
        RECT 520.1000 696.1200 522.1000 698.1200 ;
        RECT 528.2500 681.9300 530.2500 683.9300 ;
        RECT 536.4000 681.9300 538.4000 683.9300 ;
        RECT 544.5500 681.9300 546.5500 683.9300 ;
        RECT 552.7000 681.9300 554.7000 683.9300 ;
        RECT 552.7000 674.8350 554.7000 676.8350 ;
        RECT 544.5500 674.8350 546.5500 676.8350 ;
        RECT 536.4000 674.8350 538.4000 676.8350 ;
        RECT 528.2500 674.8350 530.2500 676.8350 ;
        RECT 552.7000 667.7400 554.7000 669.7400 ;
        RECT 544.5500 667.7400 546.5500 669.7400 ;
        RECT 536.4000 667.7400 538.4000 669.7400 ;
        RECT 528.2500 667.7400 530.2500 669.7400 ;
        RECT 528.2500 689.0250 530.2500 691.0250 ;
        RECT 536.4000 689.0250 538.4000 691.0250 ;
        RECT 544.5500 689.0250 546.5500 691.0250 ;
        RECT 552.7000 689.0250 554.7000 691.0250 ;
        RECT 528.2500 696.1200 530.2500 698.1200 ;
        RECT 536.4000 696.1200 538.4000 698.1200 ;
        RECT 544.5500 696.1200 546.5500 698.1200 ;
        RECT 552.7000 696.1200 554.7000 698.1200 ;
        RECT 394.0000 717.4050 396.0000 719.4050 ;
        RECT 394.0000 703.2150 396.0000 705.2150 ;
        RECT 394.0000 710.3100 396.0000 712.3100 ;
        RECT 414.1500 703.2150 416.1500 705.2150 ;
        RECT 394.0000 724.5000 396.0000 726.0000 ;
        RECT 422.3000 703.2150 424.3000 705.2150 ;
        RECT 430.4500 703.2150 432.4500 705.2150 ;
        RECT 438.6000 703.2150 440.6000 705.2150 ;
        RECT 446.7500 703.2150 448.7500 705.2150 ;
        RECT 454.9000 703.2150 456.9000 705.2150 ;
        RECT 463.0500 703.2150 465.0500 705.2150 ;
        RECT 471.2000 703.2150 473.2000 705.2150 ;
        RECT 479.3500 703.2150 481.3500 705.2150 ;
        RECT 487.5000 703.2150 489.5000 705.2150 ;
        RECT 528.2500 703.2150 530.2500 705.2150 ;
        RECT 495.6500 703.2150 497.6500 705.2150 ;
        RECT 503.8000 703.2150 505.8000 705.2150 ;
        RECT 511.9500 703.2150 513.9500 705.2150 ;
        RECT 520.1000 703.2150 522.1000 705.2150 ;
        RECT 536.4000 703.2150 538.4000 705.2150 ;
        RECT 544.5500 703.2150 546.5500 705.2150 ;
        RECT 552.7000 703.2150 554.7000 705.2150 ;
        RECT 6.0000 979.9200 8.0000 981.9200 ;
        RECT 6.0000 908.9700 8.0000 910.9700 ;
        RECT 6.0000 873.4950 8.0000 875.4950 ;
        RECT 6.0000 845.1150 8.0000 847.1150 ;
        RECT 6.0000 852.2100 8.0000 854.2100 ;
        RECT 6.0000 859.3050 8.0000 861.3050 ;
        RECT 6.0000 866.4000 8.0000 868.4000 ;
        RECT 6.0000 880.5900 8.0000 882.5900 ;
        RECT 6.0000 887.6850 8.0000 889.6850 ;
        RECT 6.0000 894.7800 8.0000 896.7800 ;
        RECT 6.0000 901.8750 8.0000 903.8750 ;
        RECT 6.0000 944.4450 8.0000 946.4450 ;
        RECT 6.0000 916.0650 8.0000 918.0650 ;
        RECT 6.0000 923.1600 8.0000 925.1600 ;
        RECT 6.0000 930.2550 8.0000 932.2550 ;
        RECT 6.0000 937.3500 8.0000 939.3500 ;
        RECT 6.0000 951.5400 8.0000 953.5400 ;
        RECT 6.0000 958.6350 8.0000 960.6350 ;
        RECT 6.0000 965.7300 8.0000 967.7300 ;
        RECT 6.0000 972.8250 8.0000 974.8250 ;
        RECT 6.0000 987.0150 8.0000 989.0150 ;
        RECT 6.0000 994.1100 8.0000 996.1100 ;
        RECT 6.0000 1001.2050 8.0000 1003.2050 ;
        RECT 6.0000 1008.3000 8.0000 1010.3000 ;
        RECT 6.0000 1022.4900 8.0000 1024.4900 ;
        RECT 6.0000 1015.3950 8.0000 1017.3950 ;
        RECT 6.0000 1029.5850 8.0000 1031.5850 ;
        RECT 6.0000 1043.7750 8.0000 1045.7750 ;
        RECT 6.0000 1036.6800 8.0000 1038.6800 ;
        RECT 6.0000 1057.9650 8.0000 1059.9650 ;
        RECT 6.0000 1050.8700 8.0000 1052.8700 ;
        RECT 6.0000 1065.0600 8.0000 1067.0600 ;
        RECT 6.0000 1072.1550 8.0000 1074.1550 ;
        RECT 6.0000 1079.2500 8.0000 1081.2500 ;
        RECT 6.0000 1100.5350 8.0000 1102.5350 ;
        RECT 6.0000 1093.4400 8.0000 1095.4400 ;
        RECT 6.0000 1086.3450 8.0000 1088.3450 ;
        RECT 6.0000 1107.6300 8.0000 1109.6300 ;
        RECT 1112.0000 838.0200 1114.0000 840.0200 ;
        RECT 699.4000 625.1700 701.4000 627.1700 ;
        RECT 699.4000 618.0750 701.4000 620.0750 ;
        RECT 699.4000 610.9800 701.4000 612.9800 ;
        RECT 699.4000 603.8850 701.4000 605.8850 ;
        RECT 699.4000 596.7900 701.4000 598.7900 ;
        RECT 699.4000 589.6950 701.4000 591.6950 ;
        RECT 699.4000 582.6000 701.4000 584.6000 ;
        RECT 699.4000 575.5050 701.4000 577.5050 ;
        RECT 699.4000 568.4100 701.4000 570.4100 ;
        RECT 699.4000 561.3150 701.4000 563.3150 ;
        RECT 699.4000 632.2650 701.4000 634.2650 ;
        RECT 699.4000 639.3600 701.4000 641.3600 ;
        RECT 699.4000 646.4550 701.4000 648.4550 ;
        RECT 699.4000 653.5500 701.4000 655.5500 ;
        RECT 699.4000 660.6450 701.4000 662.6450 ;
        RECT 699.4000 667.7400 701.4000 669.7400 ;
        RECT 699.4000 674.8350 701.4000 676.8350 ;
        RECT 699.4000 681.9300 701.4000 683.9300 ;
        RECT 699.4000 689.0250 701.4000 691.0250 ;
        RECT 699.4000 696.1200 701.4000 698.1200 ;
        RECT 593.4500 561.3150 595.4500 563.3150 ;
        RECT 593.4500 568.4100 595.4500 570.4100 ;
        RECT 593.4500 575.5050 595.4500 577.5050 ;
        RECT 593.4500 582.6000 595.4500 584.6000 ;
        RECT 593.4500 589.6950 595.4500 591.6950 ;
        RECT 560.8500 575.5050 562.8500 577.5050 ;
        RECT 569.0000 575.5050 571.0000 577.5050 ;
        RECT 577.1500 575.5050 579.1500 577.5050 ;
        RECT 585.3000 575.5050 587.3000 577.5050 ;
        RECT 585.3000 568.4100 587.3000 570.4100 ;
        RECT 577.1500 568.4100 579.1500 570.4100 ;
        RECT 569.0000 568.4100 571.0000 570.4100 ;
        RECT 560.8500 568.4100 562.8500 570.4100 ;
        RECT 585.3000 561.3150 587.3000 563.3150 ;
        RECT 577.1500 561.3150 579.1500 563.3150 ;
        RECT 569.0000 561.3150 571.0000 563.3150 ;
        RECT 560.8500 561.3150 562.8500 563.3150 ;
        RECT 560.8500 582.6000 562.8500 584.6000 ;
        RECT 569.0000 582.6000 571.0000 584.6000 ;
        RECT 577.1500 582.6000 579.1500 584.6000 ;
        RECT 585.3000 582.6000 587.3000 584.6000 ;
        RECT 560.8500 589.6950 562.8500 591.6950 ;
        RECT 569.0000 589.6950 571.0000 591.6950 ;
        RECT 577.1500 589.6950 579.1500 591.6950 ;
        RECT 585.3000 589.6950 587.3000 591.6950 ;
        RECT 601.6000 575.5050 603.6000 577.5050 ;
        RECT 609.7500 575.5050 611.7500 577.5050 ;
        RECT 617.9000 575.5050 619.9000 577.5050 ;
        RECT 626.0500 575.5050 628.0500 577.5050 ;
        RECT 626.0500 568.4100 628.0500 570.4100 ;
        RECT 617.9000 568.4100 619.9000 570.4100 ;
        RECT 609.7500 568.4100 611.7500 570.4100 ;
        RECT 601.6000 568.4100 603.6000 570.4100 ;
        RECT 626.0500 561.3150 628.0500 563.3150 ;
        RECT 617.9000 561.3150 619.9000 563.3150 ;
        RECT 609.7500 561.3150 611.7500 563.3150 ;
        RECT 601.6000 561.3150 603.6000 563.3150 ;
        RECT 601.6000 582.6000 603.6000 584.6000 ;
        RECT 609.7500 582.6000 611.7500 584.6000 ;
        RECT 617.9000 582.6000 619.9000 584.6000 ;
        RECT 626.0500 582.6000 628.0500 584.6000 ;
        RECT 601.6000 589.6950 603.6000 591.6950 ;
        RECT 609.7500 589.6950 611.7500 591.6950 ;
        RECT 617.9000 589.6950 619.9000 591.6950 ;
        RECT 626.0500 589.6950 628.0500 591.6950 ;
        RECT 593.4500 596.7900 595.4500 598.7900 ;
        RECT 593.4500 603.8850 595.4500 605.8850 ;
        RECT 593.4500 610.9800 595.4500 612.9800 ;
        RECT 593.4500 618.0750 595.4500 620.0750 ;
        RECT 593.4500 625.1700 595.4500 627.1700 ;
        RECT 560.8500 610.9800 562.8500 612.9800 ;
        RECT 569.0000 610.9800 571.0000 612.9800 ;
        RECT 577.1500 610.9800 579.1500 612.9800 ;
        RECT 585.3000 610.9800 587.3000 612.9800 ;
        RECT 585.3000 603.8850 587.3000 605.8850 ;
        RECT 577.1500 603.8850 579.1500 605.8850 ;
        RECT 569.0000 603.8850 571.0000 605.8850 ;
        RECT 560.8500 603.8850 562.8500 605.8850 ;
        RECT 585.3000 596.7900 587.3000 598.7900 ;
        RECT 577.1500 596.7900 579.1500 598.7900 ;
        RECT 569.0000 596.7900 571.0000 598.7900 ;
        RECT 560.8500 596.7900 562.8500 598.7900 ;
        RECT 560.8500 618.0750 562.8500 620.0750 ;
        RECT 569.0000 618.0750 571.0000 620.0750 ;
        RECT 577.1500 618.0750 579.1500 620.0750 ;
        RECT 585.3000 618.0750 587.3000 620.0750 ;
        RECT 560.8500 625.1700 562.8500 627.1700 ;
        RECT 569.0000 625.1700 571.0000 627.1700 ;
        RECT 577.1500 625.1700 579.1500 627.1700 ;
        RECT 585.3000 625.1700 587.3000 627.1700 ;
        RECT 601.6000 610.9800 603.6000 612.9800 ;
        RECT 609.7500 610.9800 611.7500 612.9800 ;
        RECT 617.9000 610.9800 619.9000 612.9800 ;
        RECT 626.0500 610.9800 628.0500 612.9800 ;
        RECT 626.0500 603.8850 628.0500 605.8850 ;
        RECT 617.9000 603.8850 619.9000 605.8850 ;
        RECT 609.7500 603.8850 611.7500 605.8850 ;
        RECT 601.6000 603.8850 603.6000 605.8850 ;
        RECT 626.0500 596.7900 628.0500 598.7900 ;
        RECT 617.9000 596.7900 619.9000 598.7900 ;
        RECT 609.7500 596.7900 611.7500 598.7900 ;
        RECT 601.6000 596.7900 603.6000 598.7900 ;
        RECT 601.6000 618.0750 603.6000 620.0750 ;
        RECT 609.7500 618.0750 611.7500 620.0750 ;
        RECT 617.9000 618.0750 619.9000 620.0750 ;
        RECT 626.0500 618.0750 628.0500 620.0750 ;
        RECT 601.6000 625.1700 603.6000 627.1700 ;
        RECT 609.7500 625.1700 611.7500 627.1700 ;
        RECT 617.9000 625.1700 619.9000 627.1700 ;
        RECT 626.0500 625.1700 628.0500 627.1700 ;
        RECT 634.2000 575.5050 636.2000 577.5050 ;
        RECT 642.3500 575.5050 644.3500 577.5050 ;
        RECT 650.5000 575.5050 652.5000 577.5050 ;
        RECT 658.6500 575.5050 660.6500 577.5050 ;
        RECT 658.6500 568.4100 660.6500 570.4100 ;
        RECT 650.5000 568.4100 652.5000 570.4100 ;
        RECT 642.3500 568.4100 644.3500 570.4100 ;
        RECT 634.2000 568.4100 636.2000 570.4100 ;
        RECT 658.6500 561.3150 660.6500 563.3150 ;
        RECT 650.5000 561.3150 652.5000 563.3150 ;
        RECT 642.3500 561.3150 644.3500 563.3150 ;
        RECT 634.2000 561.3150 636.2000 563.3150 ;
        RECT 634.2000 582.6000 636.2000 584.6000 ;
        RECT 642.3500 582.6000 644.3500 584.6000 ;
        RECT 650.5000 582.6000 652.5000 584.6000 ;
        RECT 658.6500 582.6000 660.6500 584.6000 ;
        RECT 634.2000 589.6950 636.2000 591.6950 ;
        RECT 642.3500 589.6950 644.3500 591.6950 ;
        RECT 650.5000 589.6950 652.5000 591.6950 ;
        RECT 658.6500 589.6950 660.6500 591.6950 ;
        RECT 666.8000 575.5050 668.8000 577.5050 ;
        RECT 674.9500 575.5050 676.9500 577.5050 ;
        RECT 683.1000 575.5050 685.1000 577.5050 ;
        RECT 691.2500 575.5050 693.2500 577.5050 ;
        RECT 691.2500 568.4100 693.2500 570.4100 ;
        RECT 683.1000 568.4100 685.1000 570.4100 ;
        RECT 674.9500 568.4100 676.9500 570.4100 ;
        RECT 666.8000 568.4100 668.8000 570.4100 ;
        RECT 691.2500 561.3150 693.2500 563.3150 ;
        RECT 683.1000 561.3150 685.1000 563.3150 ;
        RECT 674.9500 561.3150 676.9500 563.3150 ;
        RECT 666.8000 561.3150 668.8000 563.3150 ;
        RECT 666.8000 582.6000 668.8000 584.6000 ;
        RECT 674.9500 582.6000 676.9500 584.6000 ;
        RECT 683.1000 582.6000 685.1000 584.6000 ;
        RECT 691.2500 582.6000 693.2500 584.6000 ;
        RECT 666.8000 589.6950 668.8000 591.6950 ;
        RECT 674.9500 589.6950 676.9500 591.6950 ;
        RECT 683.1000 589.6950 685.1000 591.6950 ;
        RECT 691.2500 589.6950 693.2500 591.6950 ;
        RECT 634.2000 610.9800 636.2000 612.9800 ;
        RECT 642.3500 610.9800 644.3500 612.9800 ;
        RECT 650.5000 610.9800 652.5000 612.9800 ;
        RECT 658.6500 610.9800 660.6500 612.9800 ;
        RECT 658.6500 603.8850 660.6500 605.8850 ;
        RECT 650.5000 603.8850 652.5000 605.8850 ;
        RECT 642.3500 603.8850 644.3500 605.8850 ;
        RECT 634.2000 603.8850 636.2000 605.8850 ;
        RECT 658.6500 596.7900 660.6500 598.7900 ;
        RECT 650.5000 596.7900 652.5000 598.7900 ;
        RECT 642.3500 596.7900 644.3500 598.7900 ;
        RECT 634.2000 596.7900 636.2000 598.7900 ;
        RECT 634.2000 618.0750 636.2000 620.0750 ;
        RECT 642.3500 618.0750 644.3500 620.0750 ;
        RECT 650.5000 618.0750 652.5000 620.0750 ;
        RECT 658.6500 618.0750 660.6500 620.0750 ;
        RECT 634.2000 625.1700 636.2000 627.1700 ;
        RECT 642.3500 625.1700 644.3500 627.1700 ;
        RECT 650.5000 625.1700 652.5000 627.1700 ;
        RECT 658.6500 625.1700 660.6500 627.1700 ;
        RECT 666.8000 610.9800 668.8000 612.9800 ;
        RECT 674.9500 610.9800 676.9500 612.9800 ;
        RECT 683.1000 610.9800 685.1000 612.9800 ;
        RECT 691.2500 610.9800 693.2500 612.9800 ;
        RECT 691.2500 603.8850 693.2500 605.8850 ;
        RECT 683.1000 603.8850 685.1000 605.8850 ;
        RECT 674.9500 603.8850 676.9500 605.8850 ;
        RECT 666.8000 603.8850 668.8000 605.8850 ;
        RECT 691.2500 596.7900 693.2500 598.7900 ;
        RECT 683.1000 596.7900 685.1000 598.7900 ;
        RECT 674.9500 596.7900 676.9500 598.7900 ;
        RECT 666.8000 596.7900 668.8000 598.7900 ;
        RECT 666.8000 618.0750 668.8000 620.0750 ;
        RECT 674.9500 618.0750 676.9500 620.0750 ;
        RECT 683.1000 618.0750 685.1000 620.0750 ;
        RECT 691.2500 618.0750 693.2500 620.0750 ;
        RECT 666.8000 625.1700 668.8000 627.1700 ;
        RECT 674.9500 625.1700 676.9500 627.1700 ;
        RECT 683.1000 625.1700 685.1000 627.1700 ;
        RECT 691.2500 625.1700 693.2500 627.1700 ;
        RECT 593.4500 632.2650 595.4500 634.2650 ;
        RECT 593.4500 639.3600 595.4500 641.3600 ;
        RECT 593.4500 646.4550 595.4500 648.4550 ;
        RECT 593.4500 653.5500 595.4500 655.5500 ;
        RECT 593.4500 660.6450 595.4500 662.6450 ;
        RECT 560.8500 646.4550 562.8500 648.4550 ;
        RECT 569.0000 646.4550 571.0000 648.4550 ;
        RECT 577.1500 646.4550 579.1500 648.4550 ;
        RECT 585.3000 646.4550 587.3000 648.4550 ;
        RECT 585.3000 639.3600 587.3000 641.3600 ;
        RECT 577.1500 639.3600 579.1500 641.3600 ;
        RECT 569.0000 639.3600 571.0000 641.3600 ;
        RECT 560.8500 639.3600 562.8500 641.3600 ;
        RECT 585.3000 632.2650 587.3000 634.2650 ;
        RECT 577.1500 632.2650 579.1500 634.2650 ;
        RECT 569.0000 632.2650 571.0000 634.2650 ;
        RECT 560.8500 632.2650 562.8500 634.2650 ;
        RECT 560.8500 653.5500 562.8500 655.5500 ;
        RECT 569.0000 653.5500 571.0000 655.5500 ;
        RECT 577.1500 653.5500 579.1500 655.5500 ;
        RECT 585.3000 653.5500 587.3000 655.5500 ;
        RECT 560.8500 660.6450 562.8500 662.6450 ;
        RECT 569.0000 660.6450 571.0000 662.6450 ;
        RECT 577.1500 660.6450 579.1500 662.6450 ;
        RECT 585.3000 660.6450 587.3000 662.6450 ;
        RECT 601.6000 646.4550 603.6000 648.4550 ;
        RECT 609.7500 646.4550 611.7500 648.4550 ;
        RECT 617.9000 646.4550 619.9000 648.4550 ;
        RECT 626.0500 646.4550 628.0500 648.4550 ;
        RECT 626.0500 639.3600 628.0500 641.3600 ;
        RECT 617.9000 639.3600 619.9000 641.3600 ;
        RECT 609.7500 639.3600 611.7500 641.3600 ;
        RECT 601.6000 639.3600 603.6000 641.3600 ;
        RECT 626.0500 632.2650 628.0500 634.2650 ;
        RECT 617.9000 632.2650 619.9000 634.2650 ;
        RECT 609.7500 632.2650 611.7500 634.2650 ;
        RECT 601.6000 632.2650 603.6000 634.2650 ;
        RECT 601.6000 653.5500 603.6000 655.5500 ;
        RECT 609.7500 653.5500 611.7500 655.5500 ;
        RECT 617.9000 653.5500 619.9000 655.5500 ;
        RECT 626.0500 653.5500 628.0500 655.5500 ;
        RECT 601.6000 660.6450 603.6000 662.6450 ;
        RECT 609.7500 660.6450 611.7500 662.6450 ;
        RECT 617.9000 660.6450 619.9000 662.6450 ;
        RECT 626.0500 660.6450 628.0500 662.6450 ;
        RECT 593.4500 667.7400 595.4500 669.7400 ;
        RECT 593.4500 674.8350 595.4500 676.8350 ;
        RECT 593.4500 681.9300 595.4500 683.9300 ;
        RECT 593.4500 689.0250 595.4500 691.0250 ;
        RECT 593.4500 696.1200 595.4500 698.1200 ;
        RECT 560.8500 681.9300 562.8500 683.9300 ;
        RECT 569.0000 681.9300 571.0000 683.9300 ;
        RECT 577.1500 681.9300 579.1500 683.9300 ;
        RECT 585.3000 681.9300 587.3000 683.9300 ;
        RECT 585.3000 674.8350 587.3000 676.8350 ;
        RECT 577.1500 674.8350 579.1500 676.8350 ;
        RECT 569.0000 674.8350 571.0000 676.8350 ;
        RECT 560.8500 674.8350 562.8500 676.8350 ;
        RECT 585.3000 667.7400 587.3000 669.7400 ;
        RECT 577.1500 667.7400 579.1500 669.7400 ;
        RECT 569.0000 667.7400 571.0000 669.7400 ;
        RECT 560.8500 667.7400 562.8500 669.7400 ;
        RECT 560.8500 689.0250 562.8500 691.0250 ;
        RECT 569.0000 689.0250 571.0000 691.0250 ;
        RECT 577.1500 689.0250 579.1500 691.0250 ;
        RECT 585.3000 689.0250 587.3000 691.0250 ;
        RECT 560.8500 696.1200 562.8500 698.1200 ;
        RECT 569.0000 696.1200 571.0000 698.1200 ;
        RECT 577.1500 696.1200 579.1500 698.1200 ;
        RECT 585.3000 696.1200 587.3000 698.1200 ;
        RECT 601.6000 681.9300 603.6000 683.9300 ;
        RECT 609.7500 681.9300 611.7500 683.9300 ;
        RECT 617.9000 681.9300 619.9000 683.9300 ;
        RECT 626.0500 681.9300 628.0500 683.9300 ;
        RECT 626.0500 674.8350 628.0500 676.8350 ;
        RECT 617.9000 674.8350 619.9000 676.8350 ;
        RECT 609.7500 674.8350 611.7500 676.8350 ;
        RECT 601.6000 674.8350 603.6000 676.8350 ;
        RECT 626.0500 667.7400 628.0500 669.7400 ;
        RECT 617.9000 667.7400 619.9000 669.7400 ;
        RECT 609.7500 667.7400 611.7500 669.7400 ;
        RECT 601.6000 667.7400 603.6000 669.7400 ;
        RECT 601.6000 689.0250 603.6000 691.0250 ;
        RECT 609.7500 689.0250 611.7500 691.0250 ;
        RECT 617.9000 689.0250 619.9000 691.0250 ;
        RECT 626.0500 689.0250 628.0500 691.0250 ;
        RECT 601.6000 696.1200 603.6000 698.1200 ;
        RECT 609.7500 696.1200 611.7500 698.1200 ;
        RECT 617.9000 696.1200 619.9000 698.1200 ;
        RECT 626.0500 696.1200 628.0500 698.1200 ;
        RECT 634.2000 646.4550 636.2000 648.4550 ;
        RECT 642.3500 646.4550 644.3500 648.4550 ;
        RECT 650.5000 646.4550 652.5000 648.4550 ;
        RECT 658.6500 646.4550 660.6500 648.4550 ;
        RECT 658.6500 639.3600 660.6500 641.3600 ;
        RECT 650.5000 639.3600 652.5000 641.3600 ;
        RECT 642.3500 639.3600 644.3500 641.3600 ;
        RECT 634.2000 639.3600 636.2000 641.3600 ;
        RECT 658.6500 632.2650 660.6500 634.2650 ;
        RECT 650.5000 632.2650 652.5000 634.2650 ;
        RECT 642.3500 632.2650 644.3500 634.2650 ;
        RECT 634.2000 632.2650 636.2000 634.2650 ;
        RECT 634.2000 653.5500 636.2000 655.5500 ;
        RECT 642.3500 653.5500 644.3500 655.5500 ;
        RECT 650.5000 653.5500 652.5000 655.5500 ;
        RECT 658.6500 653.5500 660.6500 655.5500 ;
        RECT 634.2000 660.6450 636.2000 662.6450 ;
        RECT 642.3500 660.6450 644.3500 662.6450 ;
        RECT 650.5000 660.6450 652.5000 662.6450 ;
        RECT 658.6500 660.6450 660.6500 662.6450 ;
        RECT 666.8000 646.4550 668.8000 648.4550 ;
        RECT 674.9500 646.4550 676.9500 648.4550 ;
        RECT 683.1000 646.4550 685.1000 648.4550 ;
        RECT 691.2500 646.4550 693.2500 648.4550 ;
        RECT 691.2500 639.3600 693.2500 641.3600 ;
        RECT 683.1000 639.3600 685.1000 641.3600 ;
        RECT 674.9500 639.3600 676.9500 641.3600 ;
        RECT 666.8000 639.3600 668.8000 641.3600 ;
        RECT 691.2500 632.2650 693.2500 634.2650 ;
        RECT 683.1000 632.2650 685.1000 634.2650 ;
        RECT 674.9500 632.2650 676.9500 634.2650 ;
        RECT 666.8000 632.2650 668.8000 634.2650 ;
        RECT 666.8000 653.5500 668.8000 655.5500 ;
        RECT 674.9500 653.5500 676.9500 655.5500 ;
        RECT 683.1000 653.5500 685.1000 655.5500 ;
        RECT 691.2500 653.5500 693.2500 655.5500 ;
        RECT 666.8000 660.6450 668.8000 662.6450 ;
        RECT 674.9500 660.6450 676.9500 662.6450 ;
        RECT 683.1000 660.6450 685.1000 662.6450 ;
        RECT 691.2500 660.6450 693.2500 662.6450 ;
        RECT 634.2000 681.9300 636.2000 683.9300 ;
        RECT 642.3500 681.9300 644.3500 683.9300 ;
        RECT 650.5000 681.9300 652.5000 683.9300 ;
        RECT 658.6500 681.9300 660.6500 683.9300 ;
        RECT 658.6500 674.8350 660.6500 676.8350 ;
        RECT 650.5000 674.8350 652.5000 676.8350 ;
        RECT 642.3500 674.8350 644.3500 676.8350 ;
        RECT 634.2000 674.8350 636.2000 676.8350 ;
        RECT 658.6500 667.7400 660.6500 669.7400 ;
        RECT 650.5000 667.7400 652.5000 669.7400 ;
        RECT 642.3500 667.7400 644.3500 669.7400 ;
        RECT 634.2000 667.7400 636.2000 669.7400 ;
        RECT 634.2000 689.0250 636.2000 691.0250 ;
        RECT 642.3500 689.0250 644.3500 691.0250 ;
        RECT 650.5000 689.0250 652.5000 691.0250 ;
        RECT 658.6500 689.0250 660.6500 691.0250 ;
        RECT 634.2000 696.1200 636.2000 698.1200 ;
        RECT 642.3500 696.1200 644.3500 698.1200 ;
        RECT 650.5000 696.1200 652.5000 698.1200 ;
        RECT 658.6500 696.1200 660.6500 698.1200 ;
        RECT 666.8000 681.9300 668.8000 683.9300 ;
        RECT 674.9500 681.9300 676.9500 683.9300 ;
        RECT 683.1000 681.9300 685.1000 683.9300 ;
        RECT 691.2500 681.9300 693.2500 683.9300 ;
        RECT 691.2500 674.8350 693.2500 676.8350 ;
        RECT 683.1000 674.8350 685.1000 676.8350 ;
        RECT 674.9500 674.8350 676.9500 676.8350 ;
        RECT 666.8000 674.8350 668.8000 676.8350 ;
        RECT 691.2500 667.7400 693.2500 669.7400 ;
        RECT 683.1000 667.7400 685.1000 669.7400 ;
        RECT 674.9500 667.7400 676.9500 669.7400 ;
        RECT 666.8000 667.7400 668.8000 669.7400 ;
        RECT 666.8000 689.0250 668.8000 691.0250 ;
        RECT 674.9500 689.0250 676.9500 691.0250 ;
        RECT 683.1000 689.0250 685.1000 691.0250 ;
        RECT 691.2500 689.0250 693.2500 691.0250 ;
        RECT 666.8000 696.1200 668.8000 698.1200 ;
        RECT 674.9500 696.1200 676.9500 698.1200 ;
        RECT 683.1000 696.1200 685.1000 698.1200 ;
        RECT 691.2500 696.1200 693.2500 698.1200 ;
        RECT 707.5500 575.5050 709.5500 577.5050 ;
        RECT 715.7000 575.5050 717.7000 577.5050 ;
        RECT 723.8500 575.5050 725.8500 577.5050 ;
        RECT 732.0000 575.5050 734.0000 577.5050 ;
        RECT 732.0000 568.4100 734.0000 570.4100 ;
        RECT 723.8500 568.4100 725.8500 570.4100 ;
        RECT 715.7000 568.4100 717.7000 570.4100 ;
        RECT 707.5500 568.4100 709.5500 570.4100 ;
        RECT 732.0000 561.3150 734.0000 563.3150 ;
        RECT 723.8500 561.3150 725.8500 563.3150 ;
        RECT 715.7000 561.3150 717.7000 563.3150 ;
        RECT 707.5500 561.3150 709.5500 563.3150 ;
        RECT 707.5500 582.6000 709.5500 584.6000 ;
        RECT 715.7000 582.6000 717.7000 584.6000 ;
        RECT 723.8500 582.6000 725.8500 584.6000 ;
        RECT 732.0000 582.6000 734.0000 584.6000 ;
        RECT 707.5500 589.6950 709.5500 591.6950 ;
        RECT 715.7000 589.6950 717.7000 591.6950 ;
        RECT 723.8500 589.6950 725.8500 591.6950 ;
        RECT 732.0000 589.6950 734.0000 591.6950 ;
        RECT 740.1500 575.5050 742.1500 577.5050 ;
        RECT 748.3000 575.5050 750.3000 577.5050 ;
        RECT 756.4500 575.5050 758.4500 577.5050 ;
        RECT 764.6000 575.5050 766.6000 577.5050 ;
        RECT 764.6000 568.4100 766.6000 570.4100 ;
        RECT 756.4500 568.4100 758.4500 570.4100 ;
        RECT 748.3000 568.4100 750.3000 570.4100 ;
        RECT 740.1500 568.4100 742.1500 570.4100 ;
        RECT 764.6000 561.3150 766.6000 563.3150 ;
        RECT 756.4500 561.3150 758.4500 563.3150 ;
        RECT 748.3000 561.3150 750.3000 563.3150 ;
        RECT 740.1500 561.3150 742.1500 563.3150 ;
        RECT 740.1500 582.6000 742.1500 584.6000 ;
        RECT 748.3000 582.6000 750.3000 584.6000 ;
        RECT 756.4500 582.6000 758.4500 584.6000 ;
        RECT 764.6000 582.6000 766.6000 584.6000 ;
        RECT 740.1500 589.6950 742.1500 591.6950 ;
        RECT 748.3000 589.6950 750.3000 591.6950 ;
        RECT 756.4500 589.6950 758.4500 591.6950 ;
        RECT 764.6000 589.6950 766.6000 591.6950 ;
        RECT 707.5500 610.9800 709.5500 612.9800 ;
        RECT 715.7000 610.9800 717.7000 612.9800 ;
        RECT 723.8500 610.9800 725.8500 612.9800 ;
        RECT 732.0000 610.9800 734.0000 612.9800 ;
        RECT 732.0000 603.8850 734.0000 605.8850 ;
        RECT 723.8500 603.8850 725.8500 605.8850 ;
        RECT 715.7000 603.8850 717.7000 605.8850 ;
        RECT 707.5500 603.8850 709.5500 605.8850 ;
        RECT 732.0000 596.7900 734.0000 598.7900 ;
        RECT 723.8500 596.7900 725.8500 598.7900 ;
        RECT 715.7000 596.7900 717.7000 598.7900 ;
        RECT 707.5500 596.7900 709.5500 598.7900 ;
        RECT 707.5500 618.0750 709.5500 620.0750 ;
        RECT 715.7000 618.0750 717.7000 620.0750 ;
        RECT 723.8500 618.0750 725.8500 620.0750 ;
        RECT 732.0000 618.0750 734.0000 620.0750 ;
        RECT 707.5500 625.1700 709.5500 627.1700 ;
        RECT 715.7000 625.1700 717.7000 627.1700 ;
        RECT 723.8500 625.1700 725.8500 627.1700 ;
        RECT 732.0000 625.1700 734.0000 627.1700 ;
        RECT 740.1500 610.9800 742.1500 612.9800 ;
        RECT 748.3000 610.9800 750.3000 612.9800 ;
        RECT 756.4500 610.9800 758.4500 612.9800 ;
        RECT 764.6000 610.9800 766.6000 612.9800 ;
        RECT 764.6000 603.8850 766.6000 605.8850 ;
        RECT 756.4500 603.8850 758.4500 605.8850 ;
        RECT 748.3000 603.8850 750.3000 605.8850 ;
        RECT 740.1500 603.8850 742.1500 605.8850 ;
        RECT 764.6000 596.7900 766.6000 598.7900 ;
        RECT 756.4500 596.7900 758.4500 598.7900 ;
        RECT 748.3000 596.7900 750.3000 598.7900 ;
        RECT 740.1500 596.7900 742.1500 598.7900 ;
        RECT 740.1500 618.0750 742.1500 620.0750 ;
        RECT 748.3000 618.0750 750.3000 620.0750 ;
        RECT 756.4500 618.0750 758.4500 620.0750 ;
        RECT 764.6000 618.0750 766.6000 620.0750 ;
        RECT 740.1500 625.1700 742.1500 627.1700 ;
        RECT 748.3000 625.1700 750.3000 627.1700 ;
        RECT 756.4500 625.1700 758.4500 627.1700 ;
        RECT 764.6000 625.1700 766.6000 627.1700 ;
        RECT 772.7500 575.5050 774.7500 577.5050 ;
        RECT 780.9000 575.5050 782.9000 577.5050 ;
        RECT 789.0500 575.5050 791.0500 577.5050 ;
        RECT 797.2000 575.5050 799.2000 577.5050 ;
        RECT 797.2000 568.4100 799.2000 570.4100 ;
        RECT 789.0500 568.4100 791.0500 570.4100 ;
        RECT 780.9000 568.4100 782.9000 570.4100 ;
        RECT 772.7500 568.4100 774.7500 570.4100 ;
        RECT 797.2000 561.3150 799.2000 563.3150 ;
        RECT 789.0500 561.3150 791.0500 563.3150 ;
        RECT 780.9000 561.3150 782.9000 563.3150 ;
        RECT 772.7500 561.3150 774.7500 563.3150 ;
        RECT 772.7500 582.6000 774.7500 584.6000 ;
        RECT 780.9000 582.6000 782.9000 584.6000 ;
        RECT 789.0500 582.6000 791.0500 584.6000 ;
        RECT 797.2000 582.6000 799.2000 584.6000 ;
        RECT 772.7500 589.6950 774.7500 591.6950 ;
        RECT 780.9000 589.6950 782.9000 591.6950 ;
        RECT 789.0500 589.6950 791.0500 591.6950 ;
        RECT 797.2000 589.6950 799.2000 591.6950 ;
        RECT 805.3500 575.5050 807.3500 577.5050 ;
        RECT 813.5000 575.5050 815.5000 577.5050 ;
        RECT 821.6500 575.5050 823.6500 577.5050 ;
        RECT 829.8000 575.5050 831.8000 577.5050 ;
        RECT 837.9500 575.5050 839.9500 577.5050 ;
        RECT 837.9500 561.3150 839.9500 563.3150 ;
        RECT 829.8000 561.3150 831.8000 563.3150 ;
        RECT 821.6500 561.3150 823.6500 563.3150 ;
        RECT 813.5000 561.3150 815.5000 563.3150 ;
        RECT 805.3500 561.3150 807.3500 563.3150 ;
        RECT 805.3500 568.4100 807.3500 570.4100 ;
        RECT 813.5000 568.4100 815.5000 570.4100 ;
        RECT 821.6500 568.4100 823.6500 570.4100 ;
        RECT 829.8000 568.4100 831.8000 570.4100 ;
        RECT 837.9500 568.4100 839.9500 570.4100 ;
        RECT 805.3500 582.6000 807.3500 584.6000 ;
        RECT 813.5000 582.6000 815.5000 584.6000 ;
        RECT 821.6500 582.6000 823.6500 584.6000 ;
        RECT 829.8000 582.6000 831.8000 584.6000 ;
        RECT 837.9500 582.6000 839.9500 584.6000 ;
        RECT 805.3500 589.6950 807.3500 591.6950 ;
        RECT 813.5000 589.6950 815.5000 591.6950 ;
        RECT 821.6500 589.6950 823.6500 591.6950 ;
        RECT 829.8000 589.6950 831.8000 591.6950 ;
        RECT 837.9500 589.6950 839.9500 591.6950 ;
        RECT 772.7500 610.9800 774.7500 612.9800 ;
        RECT 780.9000 610.9800 782.9000 612.9800 ;
        RECT 789.0500 610.9800 791.0500 612.9800 ;
        RECT 797.2000 610.9800 799.2000 612.9800 ;
        RECT 797.2000 603.8850 799.2000 605.8850 ;
        RECT 789.0500 603.8850 791.0500 605.8850 ;
        RECT 780.9000 603.8850 782.9000 605.8850 ;
        RECT 772.7500 603.8850 774.7500 605.8850 ;
        RECT 797.2000 596.7900 799.2000 598.7900 ;
        RECT 789.0500 596.7900 791.0500 598.7900 ;
        RECT 780.9000 596.7900 782.9000 598.7900 ;
        RECT 772.7500 596.7900 774.7500 598.7900 ;
        RECT 772.7500 618.0750 774.7500 620.0750 ;
        RECT 780.9000 618.0750 782.9000 620.0750 ;
        RECT 789.0500 618.0750 791.0500 620.0750 ;
        RECT 797.2000 618.0750 799.2000 620.0750 ;
        RECT 772.7500 625.1700 774.7500 627.1700 ;
        RECT 780.9000 625.1700 782.9000 627.1700 ;
        RECT 789.0500 625.1700 791.0500 627.1700 ;
        RECT 797.2000 625.1700 799.2000 627.1700 ;
        RECT 805.3500 610.9800 807.3500 612.9800 ;
        RECT 813.5000 610.9800 815.5000 612.9800 ;
        RECT 821.6500 610.9800 823.6500 612.9800 ;
        RECT 829.8000 610.9800 831.8000 612.9800 ;
        RECT 837.9500 610.9800 839.9500 612.9800 ;
        RECT 837.9500 596.7900 839.9500 598.7900 ;
        RECT 829.8000 596.7900 831.8000 598.7900 ;
        RECT 821.6500 596.7900 823.6500 598.7900 ;
        RECT 813.5000 596.7900 815.5000 598.7900 ;
        RECT 805.3500 596.7900 807.3500 598.7900 ;
        RECT 805.3500 603.8850 807.3500 605.8850 ;
        RECT 813.5000 603.8850 815.5000 605.8850 ;
        RECT 821.6500 603.8850 823.6500 605.8850 ;
        RECT 829.8000 603.8850 831.8000 605.8850 ;
        RECT 837.9500 603.8850 839.9500 605.8850 ;
        RECT 805.3500 618.0750 807.3500 620.0750 ;
        RECT 813.5000 618.0750 815.5000 620.0750 ;
        RECT 821.6500 618.0750 823.6500 620.0750 ;
        RECT 829.8000 618.0750 831.8000 620.0750 ;
        RECT 837.9500 618.0750 839.9500 620.0750 ;
        RECT 805.3500 625.1700 807.3500 627.1700 ;
        RECT 813.5000 625.1700 815.5000 627.1700 ;
        RECT 821.6500 625.1700 823.6500 627.1700 ;
        RECT 829.8000 625.1700 831.8000 627.1700 ;
        RECT 837.9500 625.1700 839.9500 627.1700 ;
        RECT 707.5500 646.4550 709.5500 648.4550 ;
        RECT 715.7000 646.4550 717.7000 648.4550 ;
        RECT 723.8500 646.4550 725.8500 648.4550 ;
        RECT 732.0000 646.4550 734.0000 648.4550 ;
        RECT 732.0000 639.3600 734.0000 641.3600 ;
        RECT 723.8500 639.3600 725.8500 641.3600 ;
        RECT 715.7000 639.3600 717.7000 641.3600 ;
        RECT 707.5500 639.3600 709.5500 641.3600 ;
        RECT 732.0000 632.2650 734.0000 634.2650 ;
        RECT 723.8500 632.2650 725.8500 634.2650 ;
        RECT 715.7000 632.2650 717.7000 634.2650 ;
        RECT 707.5500 632.2650 709.5500 634.2650 ;
        RECT 707.5500 653.5500 709.5500 655.5500 ;
        RECT 715.7000 653.5500 717.7000 655.5500 ;
        RECT 723.8500 653.5500 725.8500 655.5500 ;
        RECT 732.0000 653.5500 734.0000 655.5500 ;
        RECT 707.5500 660.6450 709.5500 662.6450 ;
        RECT 715.7000 660.6450 717.7000 662.6450 ;
        RECT 723.8500 660.6450 725.8500 662.6450 ;
        RECT 732.0000 660.6450 734.0000 662.6450 ;
        RECT 740.1500 646.4550 742.1500 648.4550 ;
        RECT 748.3000 646.4550 750.3000 648.4550 ;
        RECT 756.4500 646.4550 758.4500 648.4550 ;
        RECT 764.6000 646.4550 766.6000 648.4550 ;
        RECT 764.6000 639.3600 766.6000 641.3600 ;
        RECT 756.4500 639.3600 758.4500 641.3600 ;
        RECT 748.3000 639.3600 750.3000 641.3600 ;
        RECT 740.1500 639.3600 742.1500 641.3600 ;
        RECT 764.6000 632.2650 766.6000 634.2650 ;
        RECT 756.4500 632.2650 758.4500 634.2650 ;
        RECT 748.3000 632.2650 750.3000 634.2650 ;
        RECT 740.1500 632.2650 742.1500 634.2650 ;
        RECT 740.1500 653.5500 742.1500 655.5500 ;
        RECT 748.3000 653.5500 750.3000 655.5500 ;
        RECT 756.4500 653.5500 758.4500 655.5500 ;
        RECT 764.6000 653.5500 766.6000 655.5500 ;
        RECT 740.1500 660.6450 742.1500 662.6450 ;
        RECT 748.3000 660.6450 750.3000 662.6450 ;
        RECT 756.4500 660.6450 758.4500 662.6450 ;
        RECT 764.6000 660.6450 766.6000 662.6450 ;
        RECT 707.5500 681.9300 709.5500 683.9300 ;
        RECT 715.7000 681.9300 717.7000 683.9300 ;
        RECT 723.8500 681.9300 725.8500 683.9300 ;
        RECT 732.0000 681.9300 734.0000 683.9300 ;
        RECT 732.0000 674.8350 734.0000 676.8350 ;
        RECT 723.8500 674.8350 725.8500 676.8350 ;
        RECT 715.7000 674.8350 717.7000 676.8350 ;
        RECT 707.5500 674.8350 709.5500 676.8350 ;
        RECT 732.0000 667.7400 734.0000 669.7400 ;
        RECT 723.8500 667.7400 725.8500 669.7400 ;
        RECT 715.7000 667.7400 717.7000 669.7400 ;
        RECT 707.5500 667.7400 709.5500 669.7400 ;
        RECT 707.5500 689.0250 709.5500 691.0250 ;
        RECT 715.7000 689.0250 717.7000 691.0250 ;
        RECT 723.8500 689.0250 725.8500 691.0250 ;
        RECT 732.0000 689.0250 734.0000 691.0250 ;
        RECT 707.5500 696.1200 709.5500 698.1200 ;
        RECT 715.7000 696.1200 717.7000 698.1200 ;
        RECT 723.8500 696.1200 725.8500 698.1200 ;
        RECT 732.0000 696.1200 734.0000 698.1200 ;
        RECT 740.1500 681.9300 742.1500 683.9300 ;
        RECT 748.3000 681.9300 750.3000 683.9300 ;
        RECT 756.4500 681.9300 758.4500 683.9300 ;
        RECT 764.6000 681.9300 766.6000 683.9300 ;
        RECT 764.6000 674.8350 766.6000 676.8350 ;
        RECT 756.4500 674.8350 758.4500 676.8350 ;
        RECT 748.3000 674.8350 750.3000 676.8350 ;
        RECT 740.1500 674.8350 742.1500 676.8350 ;
        RECT 764.6000 667.7400 766.6000 669.7400 ;
        RECT 756.4500 667.7400 758.4500 669.7400 ;
        RECT 748.3000 667.7400 750.3000 669.7400 ;
        RECT 740.1500 667.7400 742.1500 669.7400 ;
        RECT 740.1500 689.0250 742.1500 691.0250 ;
        RECT 748.3000 689.0250 750.3000 691.0250 ;
        RECT 756.4500 689.0250 758.4500 691.0250 ;
        RECT 764.6000 689.0250 766.6000 691.0250 ;
        RECT 740.1500 696.1200 742.1500 698.1200 ;
        RECT 748.3000 696.1200 750.3000 698.1200 ;
        RECT 756.4500 696.1200 758.4500 698.1200 ;
        RECT 764.6000 696.1200 766.6000 698.1200 ;
        RECT 772.7500 646.4550 774.7500 648.4550 ;
        RECT 780.9000 646.4550 782.9000 648.4550 ;
        RECT 789.0500 646.4550 791.0500 648.4550 ;
        RECT 797.2000 646.4550 799.2000 648.4550 ;
        RECT 797.2000 639.3600 799.2000 641.3600 ;
        RECT 789.0500 639.3600 791.0500 641.3600 ;
        RECT 780.9000 639.3600 782.9000 641.3600 ;
        RECT 772.7500 639.3600 774.7500 641.3600 ;
        RECT 797.2000 632.2650 799.2000 634.2650 ;
        RECT 789.0500 632.2650 791.0500 634.2650 ;
        RECT 780.9000 632.2650 782.9000 634.2650 ;
        RECT 772.7500 632.2650 774.7500 634.2650 ;
        RECT 772.7500 653.5500 774.7500 655.5500 ;
        RECT 780.9000 653.5500 782.9000 655.5500 ;
        RECT 789.0500 653.5500 791.0500 655.5500 ;
        RECT 797.2000 653.5500 799.2000 655.5500 ;
        RECT 772.7500 660.6450 774.7500 662.6450 ;
        RECT 780.9000 660.6450 782.9000 662.6450 ;
        RECT 789.0500 660.6450 791.0500 662.6450 ;
        RECT 797.2000 660.6450 799.2000 662.6450 ;
        RECT 805.3500 646.4550 807.3500 648.4550 ;
        RECT 813.5000 646.4550 815.5000 648.4550 ;
        RECT 821.6500 646.4550 823.6500 648.4550 ;
        RECT 829.8000 646.4550 831.8000 648.4550 ;
        RECT 837.9500 646.4550 839.9500 648.4550 ;
        RECT 837.9500 632.2650 839.9500 634.2650 ;
        RECT 829.8000 632.2650 831.8000 634.2650 ;
        RECT 821.6500 632.2650 823.6500 634.2650 ;
        RECT 813.5000 632.2650 815.5000 634.2650 ;
        RECT 805.3500 632.2650 807.3500 634.2650 ;
        RECT 805.3500 639.3600 807.3500 641.3600 ;
        RECT 813.5000 639.3600 815.5000 641.3600 ;
        RECT 821.6500 639.3600 823.6500 641.3600 ;
        RECT 829.8000 639.3600 831.8000 641.3600 ;
        RECT 837.9500 639.3600 839.9500 641.3600 ;
        RECT 805.3500 653.5500 807.3500 655.5500 ;
        RECT 813.5000 653.5500 815.5000 655.5500 ;
        RECT 821.6500 653.5500 823.6500 655.5500 ;
        RECT 829.8000 653.5500 831.8000 655.5500 ;
        RECT 837.9500 653.5500 839.9500 655.5500 ;
        RECT 805.3500 660.6450 807.3500 662.6450 ;
        RECT 813.5000 660.6450 815.5000 662.6450 ;
        RECT 821.6500 660.6450 823.6500 662.6450 ;
        RECT 829.8000 660.6450 831.8000 662.6450 ;
        RECT 837.9500 660.6450 839.9500 662.6450 ;
        RECT 772.7500 681.9300 774.7500 683.9300 ;
        RECT 780.9000 681.9300 782.9000 683.9300 ;
        RECT 789.0500 681.9300 791.0500 683.9300 ;
        RECT 797.2000 681.9300 799.2000 683.9300 ;
        RECT 797.2000 674.8350 799.2000 676.8350 ;
        RECT 789.0500 674.8350 791.0500 676.8350 ;
        RECT 780.9000 674.8350 782.9000 676.8350 ;
        RECT 772.7500 674.8350 774.7500 676.8350 ;
        RECT 797.2000 667.7400 799.2000 669.7400 ;
        RECT 789.0500 667.7400 791.0500 669.7400 ;
        RECT 780.9000 667.7400 782.9000 669.7400 ;
        RECT 772.7500 667.7400 774.7500 669.7400 ;
        RECT 772.7500 689.0250 774.7500 691.0250 ;
        RECT 780.9000 689.0250 782.9000 691.0250 ;
        RECT 789.0500 689.0250 791.0500 691.0250 ;
        RECT 797.2000 689.0250 799.2000 691.0250 ;
        RECT 772.7500 696.1200 774.7500 698.1200 ;
        RECT 780.9000 696.1200 782.9000 698.1200 ;
        RECT 789.0500 696.1200 791.0500 698.1200 ;
        RECT 797.2000 696.1200 799.2000 698.1200 ;
        RECT 805.3500 681.9300 807.3500 683.9300 ;
        RECT 813.5000 681.9300 815.5000 683.9300 ;
        RECT 821.6500 681.9300 823.6500 683.9300 ;
        RECT 829.8000 681.9300 831.8000 683.9300 ;
        RECT 837.9500 681.9300 839.9500 683.9300 ;
        RECT 837.9500 667.7400 839.9500 669.7400 ;
        RECT 829.8000 667.7400 831.8000 669.7400 ;
        RECT 821.6500 667.7400 823.6500 669.7400 ;
        RECT 813.5000 667.7400 815.5000 669.7400 ;
        RECT 805.3500 667.7400 807.3500 669.7400 ;
        RECT 805.3500 674.8350 807.3500 676.8350 ;
        RECT 813.5000 674.8350 815.5000 676.8350 ;
        RECT 821.6500 674.8350 823.6500 676.8350 ;
        RECT 829.8000 674.8350 831.8000 676.8350 ;
        RECT 837.9500 674.8350 839.9500 676.8350 ;
        RECT 805.3500 689.0250 807.3500 691.0250 ;
        RECT 813.5000 689.0250 815.5000 691.0250 ;
        RECT 821.6500 689.0250 823.6500 691.0250 ;
        RECT 829.8000 689.0250 831.8000 691.0250 ;
        RECT 837.9500 689.0250 839.9500 691.0250 ;
        RECT 805.3500 696.1200 807.3500 698.1200 ;
        RECT 813.5000 696.1200 815.5000 698.1200 ;
        RECT 821.6500 696.1200 823.6500 698.1200 ;
        RECT 829.8000 696.1200 831.8000 698.1200 ;
        RECT 837.9500 696.1200 839.9500 698.1200 ;
        RECT 699.4000 703.2150 701.4000 705.2150 ;
        RECT 560.8500 703.2150 562.8500 705.2150 ;
        RECT 569.0000 703.2150 571.0000 705.2150 ;
        RECT 577.1500 703.2150 579.1500 705.2150 ;
        RECT 585.3000 703.2150 587.3000 705.2150 ;
        RECT 593.4500 703.2150 595.4500 705.2150 ;
        RECT 601.6000 703.2150 603.6000 705.2150 ;
        RECT 609.7500 703.2150 611.7500 705.2150 ;
        RECT 617.9000 703.2150 619.9000 705.2150 ;
        RECT 626.0500 703.2150 628.0500 705.2150 ;
        RECT 666.8000 703.2150 668.8000 705.2150 ;
        RECT 634.2000 703.2150 636.2000 705.2150 ;
        RECT 642.3500 703.2150 644.3500 705.2150 ;
        RECT 650.5000 703.2150 652.5000 705.2150 ;
        RECT 658.6500 703.2150 660.6500 705.2150 ;
        RECT 674.9500 703.2150 676.9500 705.2150 ;
        RECT 683.1000 703.2150 685.1000 705.2150 ;
        RECT 691.2500 703.2150 693.2500 705.2150 ;
        RECT 707.5500 703.2150 709.5500 705.2150 ;
        RECT 715.7000 703.2150 717.7000 705.2150 ;
        RECT 723.8500 703.2150 725.8500 705.2150 ;
        RECT 732.0000 703.2150 734.0000 705.2150 ;
        RECT 740.1500 703.2150 742.1500 705.2150 ;
        RECT 748.3000 703.2150 750.3000 705.2150 ;
        RECT 756.4500 703.2150 758.4500 705.2150 ;
        RECT 764.6000 703.2150 766.6000 705.2150 ;
        RECT 813.5000 703.2150 815.5000 705.2150 ;
        RECT 772.7500 703.2150 774.7500 705.2150 ;
        RECT 780.9000 703.2150 782.9000 705.2150 ;
        RECT 789.0500 703.2150 791.0500 705.2150 ;
        RECT 797.2000 703.2150 799.2000 705.2150 ;
        RECT 805.3500 703.2150 807.3500 705.2150 ;
        RECT 821.6500 703.2150 823.6500 705.2150 ;
        RECT 829.8000 703.2150 831.8000 705.2150 ;
        RECT 837.9500 703.2150 839.9500 705.2150 ;
        RECT 846.1000 575.5050 848.1000 577.5050 ;
        RECT 854.2500 575.5050 856.2500 577.5050 ;
        RECT 862.4000 575.5050 864.4000 577.5050 ;
        RECT 870.5500 575.5050 872.5500 577.5050 ;
        RECT 870.5500 568.4100 872.5500 570.4100 ;
        RECT 862.4000 568.4100 864.4000 570.4100 ;
        RECT 854.2500 568.4100 856.2500 570.4100 ;
        RECT 846.1000 568.4100 848.1000 570.4100 ;
        RECT 870.5500 561.3150 872.5500 563.3150 ;
        RECT 862.4000 561.3150 864.4000 563.3150 ;
        RECT 854.2500 561.3150 856.2500 563.3150 ;
        RECT 846.1000 561.3150 848.1000 563.3150 ;
        RECT 846.1000 582.6000 848.1000 584.6000 ;
        RECT 854.2500 582.6000 856.2500 584.6000 ;
        RECT 862.4000 582.6000 864.4000 584.6000 ;
        RECT 870.5500 582.6000 872.5500 584.6000 ;
        RECT 846.1000 589.6950 848.1000 591.6950 ;
        RECT 854.2500 589.6950 856.2500 591.6950 ;
        RECT 862.4000 589.6950 864.4000 591.6950 ;
        RECT 870.5500 589.6950 872.5500 591.6950 ;
        RECT 878.7000 575.5050 880.7000 577.5050 ;
        RECT 886.8500 575.5050 888.8500 577.5050 ;
        RECT 895.0000 575.5050 897.0000 577.5050 ;
        RECT 903.1500 575.5050 905.1500 577.5050 ;
        RECT 903.1500 568.4100 905.1500 570.4100 ;
        RECT 895.0000 568.4100 897.0000 570.4100 ;
        RECT 886.8500 568.4100 888.8500 570.4100 ;
        RECT 878.7000 568.4100 880.7000 570.4100 ;
        RECT 903.1500 561.3150 905.1500 563.3150 ;
        RECT 895.0000 561.3150 897.0000 563.3150 ;
        RECT 886.8500 561.3150 888.8500 563.3150 ;
        RECT 878.7000 561.3150 880.7000 563.3150 ;
        RECT 878.7000 582.6000 880.7000 584.6000 ;
        RECT 886.8500 582.6000 888.8500 584.6000 ;
        RECT 895.0000 582.6000 897.0000 584.6000 ;
        RECT 903.1500 582.6000 905.1500 584.6000 ;
        RECT 878.7000 589.6950 880.7000 591.6950 ;
        RECT 886.8500 589.6950 888.8500 591.6950 ;
        RECT 895.0000 589.6950 897.0000 591.6950 ;
        RECT 903.1500 589.6950 905.1500 591.6950 ;
        RECT 846.1000 610.9800 848.1000 612.9800 ;
        RECT 854.2500 610.9800 856.2500 612.9800 ;
        RECT 862.4000 610.9800 864.4000 612.9800 ;
        RECT 870.5500 610.9800 872.5500 612.9800 ;
        RECT 870.5500 603.8850 872.5500 605.8850 ;
        RECT 862.4000 603.8850 864.4000 605.8850 ;
        RECT 854.2500 603.8850 856.2500 605.8850 ;
        RECT 846.1000 603.8850 848.1000 605.8850 ;
        RECT 870.5500 596.7900 872.5500 598.7900 ;
        RECT 862.4000 596.7900 864.4000 598.7900 ;
        RECT 854.2500 596.7900 856.2500 598.7900 ;
        RECT 846.1000 596.7900 848.1000 598.7900 ;
        RECT 846.1000 618.0750 848.1000 620.0750 ;
        RECT 854.2500 618.0750 856.2500 620.0750 ;
        RECT 862.4000 618.0750 864.4000 620.0750 ;
        RECT 870.5500 618.0750 872.5500 620.0750 ;
        RECT 846.1000 625.1700 848.1000 627.1700 ;
        RECT 854.2500 625.1700 856.2500 627.1700 ;
        RECT 862.4000 625.1700 864.4000 627.1700 ;
        RECT 870.5500 625.1700 872.5500 627.1700 ;
        RECT 878.7000 610.9800 880.7000 612.9800 ;
        RECT 886.8500 610.9800 888.8500 612.9800 ;
        RECT 895.0000 610.9800 897.0000 612.9800 ;
        RECT 903.1500 610.9800 905.1500 612.9800 ;
        RECT 903.1500 603.8850 905.1500 605.8850 ;
        RECT 895.0000 603.8850 897.0000 605.8850 ;
        RECT 886.8500 603.8850 888.8500 605.8850 ;
        RECT 878.7000 603.8850 880.7000 605.8850 ;
        RECT 903.1500 596.7900 905.1500 598.7900 ;
        RECT 895.0000 596.7900 897.0000 598.7900 ;
        RECT 886.8500 596.7900 888.8500 598.7900 ;
        RECT 878.7000 596.7900 880.7000 598.7900 ;
        RECT 878.7000 618.0750 880.7000 620.0750 ;
        RECT 886.8500 618.0750 888.8500 620.0750 ;
        RECT 895.0000 618.0750 897.0000 620.0750 ;
        RECT 903.1500 618.0750 905.1500 620.0750 ;
        RECT 878.7000 625.1700 880.7000 627.1700 ;
        RECT 886.8500 625.1700 888.8500 627.1700 ;
        RECT 895.0000 625.1700 897.0000 627.1700 ;
        RECT 903.1500 625.1700 905.1500 627.1700 ;
        RECT 943.9000 561.3150 945.9000 563.3150 ;
        RECT 943.9000 568.4100 945.9000 570.4100 ;
        RECT 943.9000 575.5050 945.9000 577.5050 ;
        RECT 943.9000 582.6000 945.9000 584.6000 ;
        RECT 943.9000 589.6950 945.9000 591.6950 ;
        RECT 911.3000 575.5050 913.3000 577.5050 ;
        RECT 919.4500 575.5050 921.4500 577.5050 ;
        RECT 927.6000 575.5050 929.6000 577.5050 ;
        RECT 935.7500 575.5050 937.7500 577.5050 ;
        RECT 935.7500 568.4100 937.7500 570.4100 ;
        RECT 927.6000 568.4100 929.6000 570.4100 ;
        RECT 919.4500 568.4100 921.4500 570.4100 ;
        RECT 911.3000 568.4100 913.3000 570.4100 ;
        RECT 935.7500 561.3150 937.7500 563.3150 ;
        RECT 927.6000 561.3150 929.6000 563.3150 ;
        RECT 919.4500 561.3150 921.4500 563.3150 ;
        RECT 911.3000 561.3150 913.3000 563.3150 ;
        RECT 911.3000 582.6000 913.3000 584.6000 ;
        RECT 919.4500 582.6000 921.4500 584.6000 ;
        RECT 927.6000 582.6000 929.6000 584.6000 ;
        RECT 935.7500 582.6000 937.7500 584.6000 ;
        RECT 911.3000 589.6950 913.3000 591.6950 ;
        RECT 919.4500 589.6950 921.4500 591.6950 ;
        RECT 927.6000 589.6950 929.6000 591.6950 ;
        RECT 935.7500 589.6950 937.7500 591.6950 ;
        RECT 952.0500 575.5050 954.0500 577.5050 ;
        RECT 960.2000 575.5050 962.2000 577.5050 ;
        RECT 968.3500 575.5050 970.3500 577.5050 ;
        RECT 976.5000 575.5050 978.5000 577.5050 ;
        RECT 976.5000 568.4100 978.5000 570.4100 ;
        RECT 968.3500 568.4100 970.3500 570.4100 ;
        RECT 960.2000 568.4100 962.2000 570.4100 ;
        RECT 952.0500 568.4100 954.0500 570.4100 ;
        RECT 976.5000 561.3150 978.5000 563.3150 ;
        RECT 968.3500 561.3150 970.3500 563.3150 ;
        RECT 960.2000 561.3150 962.2000 563.3150 ;
        RECT 952.0500 561.3150 954.0500 563.3150 ;
        RECT 952.0500 582.6000 954.0500 584.6000 ;
        RECT 960.2000 582.6000 962.2000 584.6000 ;
        RECT 968.3500 582.6000 970.3500 584.6000 ;
        RECT 976.5000 582.6000 978.5000 584.6000 ;
        RECT 952.0500 589.6950 954.0500 591.6950 ;
        RECT 960.2000 589.6950 962.2000 591.6950 ;
        RECT 968.3500 589.6950 970.3500 591.6950 ;
        RECT 976.5000 589.6950 978.5000 591.6950 ;
        RECT 943.9000 596.7900 945.9000 598.7900 ;
        RECT 943.9000 603.8850 945.9000 605.8850 ;
        RECT 943.9000 610.9800 945.9000 612.9800 ;
        RECT 943.9000 618.0750 945.9000 620.0750 ;
        RECT 943.9000 625.1700 945.9000 627.1700 ;
        RECT 911.3000 610.9800 913.3000 612.9800 ;
        RECT 919.4500 610.9800 921.4500 612.9800 ;
        RECT 927.6000 610.9800 929.6000 612.9800 ;
        RECT 935.7500 610.9800 937.7500 612.9800 ;
        RECT 935.7500 603.8850 937.7500 605.8850 ;
        RECT 927.6000 603.8850 929.6000 605.8850 ;
        RECT 919.4500 603.8850 921.4500 605.8850 ;
        RECT 911.3000 603.8850 913.3000 605.8850 ;
        RECT 935.7500 596.7900 937.7500 598.7900 ;
        RECT 927.6000 596.7900 929.6000 598.7900 ;
        RECT 919.4500 596.7900 921.4500 598.7900 ;
        RECT 911.3000 596.7900 913.3000 598.7900 ;
        RECT 911.3000 618.0750 913.3000 620.0750 ;
        RECT 919.4500 618.0750 921.4500 620.0750 ;
        RECT 927.6000 618.0750 929.6000 620.0750 ;
        RECT 935.7500 618.0750 937.7500 620.0750 ;
        RECT 911.3000 625.1700 913.3000 627.1700 ;
        RECT 919.4500 625.1700 921.4500 627.1700 ;
        RECT 927.6000 625.1700 929.6000 627.1700 ;
        RECT 935.7500 625.1700 937.7500 627.1700 ;
        RECT 952.0500 610.9800 954.0500 612.9800 ;
        RECT 960.2000 610.9800 962.2000 612.9800 ;
        RECT 968.3500 610.9800 970.3500 612.9800 ;
        RECT 976.5000 610.9800 978.5000 612.9800 ;
        RECT 976.5000 603.8850 978.5000 605.8850 ;
        RECT 968.3500 603.8850 970.3500 605.8850 ;
        RECT 960.2000 603.8850 962.2000 605.8850 ;
        RECT 952.0500 603.8850 954.0500 605.8850 ;
        RECT 976.5000 596.7900 978.5000 598.7900 ;
        RECT 968.3500 596.7900 970.3500 598.7900 ;
        RECT 960.2000 596.7900 962.2000 598.7900 ;
        RECT 952.0500 596.7900 954.0500 598.7900 ;
        RECT 952.0500 618.0750 954.0500 620.0750 ;
        RECT 960.2000 618.0750 962.2000 620.0750 ;
        RECT 968.3500 618.0750 970.3500 620.0750 ;
        RECT 976.5000 618.0750 978.5000 620.0750 ;
        RECT 952.0500 625.1700 954.0500 627.1700 ;
        RECT 960.2000 625.1700 962.2000 627.1700 ;
        RECT 968.3500 625.1700 970.3500 627.1700 ;
        RECT 976.5000 625.1700 978.5000 627.1700 ;
        RECT 846.1000 646.4550 848.1000 648.4550 ;
        RECT 854.2500 646.4550 856.2500 648.4550 ;
        RECT 862.4000 646.4550 864.4000 648.4550 ;
        RECT 870.5500 646.4550 872.5500 648.4550 ;
        RECT 870.5500 639.3600 872.5500 641.3600 ;
        RECT 862.4000 639.3600 864.4000 641.3600 ;
        RECT 854.2500 639.3600 856.2500 641.3600 ;
        RECT 846.1000 639.3600 848.1000 641.3600 ;
        RECT 870.5500 632.2650 872.5500 634.2650 ;
        RECT 862.4000 632.2650 864.4000 634.2650 ;
        RECT 854.2500 632.2650 856.2500 634.2650 ;
        RECT 846.1000 632.2650 848.1000 634.2650 ;
        RECT 846.1000 653.5500 848.1000 655.5500 ;
        RECT 854.2500 653.5500 856.2500 655.5500 ;
        RECT 862.4000 653.5500 864.4000 655.5500 ;
        RECT 870.5500 653.5500 872.5500 655.5500 ;
        RECT 846.1000 660.6450 848.1000 662.6450 ;
        RECT 854.2500 660.6450 856.2500 662.6450 ;
        RECT 862.4000 660.6450 864.4000 662.6450 ;
        RECT 870.5500 660.6450 872.5500 662.6450 ;
        RECT 878.7000 646.4550 880.7000 648.4550 ;
        RECT 886.8500 646.4550 888.8500 648.4550 ;
        RECT 895.0000 646.4550 897.0000 648.4550 ;
        RECT 903.1500 646.4550 905.1500 648.4550 ;
        RECT 903.1500 639.3600 905.1500 641.3600 ;
        RECT 895.0000 639.3600 897.0000 641.3600 ;
        RECT 886.8500 639.3600 888.8500 641.3600 ;
        RECT 878.7000 639.3600 880.7000 641.3600 ;
        RECT 903.1500 632.2650 905.1500 634.2650 ;
        RECT 895.0000 632.2650 897.0000 634.2650 ;
        RECT 886.8500 632.2650 888.8500 634.2650 ;
        RECT 878.7000 632.2650 880.7000 634.2650 ;
        RECT 878.7000 653.5500 880.7000 655.5500 ;
        RECT 886.8500 653.5500 888.8500 655.5500 ;
        RECT 895.0000 653.5500 897.0000 655.5500 ;
        RECT 903.1500 653.5500 905.1500 655.5500 ;
        RECT 878.7000 660.6450 880.7000 662.6450 ;
        RECT 886.8500 660.6450 888.8500 662.6450 ;
        RECT 895.0000 660.6450 897.0000 662.6450 ;
        RECT 903.1500 660.6450 905.1500 662.6450 ;
        RECT 846.1000 681.9300 848.1000 683.9300 ;
        RECT 854.2500 681.9300 856.2500 683.9300 ;
        RECT 862.4000 681.9300 864.4000 683.9300 ;
        RECT 870.5500 681.9300 872.5500 683.9300 ;
        RECT 870.5500 674.8350 872.5500 676.8350 ;
        RECT 862.4000 674.8350 864.4000 676.8350 ;
        RECT 854.2500 674.8350 856.2500 676.8350 ;
        RECT 846.1000 674.8350 848.1000 676.8350 ;
        RECT 870.5500 667.7400 872.5500 669.7400 ;
        RECT 862.4000 667.7400 864.4000 669.7400 ;
        RECT 854.2500 667.7400 856.2500 669.7400 ;
        RECT 846.1000 667.7400 848.1000 669.7400 ;
        RECT 846.1000 689.0250 848.1000 691.0250 ;
        RECT 854.2500 689.0250 856.2500 691.0250 ;
        RECT 862.4000 689.0250 864.4000 691.0250 ;
        RECT 870.5500 689.0250 872.5500 691.0250 ;
        RECT 846.1000 696.1200 848.1000 698.1200 ;
        RECT 854.2500 696.1200 856.2500 698.1200 ;
        RECT 862.4000 696.1200 864.4000 698.1200 ;
        RECT 870.5500 696.1200 872.5500 698.1200 ;
        RECT 878.7000 681.9300 880.7000 683.9300 ;
        RECT 886.8500 681.9300 888.8500 683.9300 ;
        RECT 895.0000 681.9300 897.0000 683.9300 ;
        RECT 903.1500 681.9300 905.1500 683.9300 ;
        RECT 903.1500 674.8350 905.1500 676.8350 ;
        RECT 895.0000 674.8350 897.0000 676.8350 ;
        RECT 886.8500 674.8350 888.8500 676.8350 ;
        RECT 878.7000 674.8350 880.7000 676.8350 ;
        RECT 903.1500 667.7400 905.1500 669.7400 ;
        RECT 895.0000 667.7400 897.0000 669.7400 ;
        RECT 886.8500 667.7400 888.8500 669.7400 ;
        RECT 878.7000 667.7400 880.7000 669.7400 ;
        RECT 878.7000 689.0250 880.7000 691.0250 ;
        RECT 886.8500 689.0250 888.8500 691.0250 ;
        RECT 895.0000 689.0250 897.0000 691.0250 ;
        RECT 903.1500 689.0250 905.1500 691.0250 ;
        RECT 878.7000 696.1200 880.7000 698.1200 ;
        RECT 886.8500 696.1200 888.8500 698.1200 ;
        RECT 895.0000 696.1200 897.0000 698.1200 ;
        RECT 903.1500 696.1200 905.1500 698.1200 ;
        RECT 943.9000 632.2650 945.9000 634.2650 ;
        RECT 943.9000 639.3600 945.9000 641.3600 ;
        RECT 943.9000 646.4550 945.9000 648.4550 ;
        RECT 943.9000 653.5500 945.9000 655.5500 ;
        RECT 943.9000 660.6450 945.9000 662.6450 ;
        RECT 911.3000 646.4550 913.3000 648.4550 ;
        RECT 919.4500 646.4550 921.4500 648.4550 ;
        RECT 927.6000 646.4550 929.6000 648.4550 ;
        RECT 935.7500 646.4550 937.7500 648.4550 ;
        RECT 935.7500 639.3600 937.7500 641.3600 ;
        RECT 927.6000 639.3600 929.6000 641.3600 ;
        RECT 919.4500 639.3600 921.4500 641.3600 ;
        RECT 911.3000 639.3600 913.3000 641.3600 ;
        RECT 935.7500 632.2650 937.7500 634.2650 ;
        RECT 927.6000 632.2650 929.6000 634.2650 ;
        RECT 919.4500 632.2650 921.4500 634.2650 ;
        RECT 911.3000 632.2650 913.3000 634.2650 ;
        RECT 911.3000 653.5500 913.3000 655.5500 ;
        RECT 919.4500 653.5500 921.4500 655.5500 ;
        RECT 927.6000 653.5500 929.6000 655.5500 ;
        RECT 935.7500 653.5500 937.7500 655.5500 ;
        RECT 911.3000 660.6450 913.3000 662.6450 ;
        RECT 919.4500 660.6450 921.4500 662.6450 ;
        RECT 927.6000 660.6450 929.6000 662.6450 ;
        RECT 935.7500 660.6450 937.7500 662.6450 ;
        RECT 952.0500 646.4550 954.0500 648.4550 ;
        RECT 960.2000 646.4550 962.2000 648.4550 ;
        RECT 968.3500 646.4550 970.3500 648.4550 ;
        RECT 976.5000 646.4550 978.5000 648.4550 ;
        RECT 976.5000 639.3600 978.5000 641.3600 ;
        RECT 968.3500 639.3600 970.3500 641.3600 ;
        RECT 960.2000 639.3600 962.2000 641.3600 ;
        RECT 952.0500 639.3600 954.0500 641.3600 ;
        RECT 976.5000 632.2650 978.5000 634.2650 ;
        RECT 968.3500 632.2650 970.3500 634.2650 ;
        RECT 960.2000 632.2650 962.2000 634.2650 ;
        RECT 952.0500 632.2650 954.0500 634.2650 ;
        RECT 952.0500 653.5500 954.0500 655.5500 ;
        RECT 960.2000 653.5500 962.2000 655.5500 ;
        RECT 968.3500 653.5500 970.3500 655.5500 ;
        RECT 976.5000 653.5500 978.5000 655.5500 ;
        RECT 952.0500 660.6450 954.0500 662.6450 ;
        RECT 960.2000 660.6450 962.2000 662.6450 ;
        RECT 968.3500 660.6450 970.3500 662.6450 ;
        RECT 976.5000 660.6450 978.5000 662.6450 ;
        RECT 943.9000 667.7400 945.9000 669.7400 ;
        RECT 943.9000 674.8350 945.9000 676.8350 ;
        RECT 943.9000 681.9300 945.9000 683.9300 ;
        RECT 943.9000 689.0250 945.9000 691.0250 ;
        RECT 943.9000 696.1200 945.9000 698.1200 ;
        RECT 911.3000 681.9300 913.3000 683.9300 ;
        RECT 919.4500 681.9300 921.4500 683.9300 ;
        RECT 927.6000 681.9300 929.6000 683.9300 ;
        RECT 935.7500 681.9300 937.7500 683.9300 ;
        RECT 935.7500 674.8350 937.7500 676.8350 ;
        RECT 927.6000 674.8350 929.6000 676.8350 ;
        RECT 919.4500 674.8350 921.4500 676.8350 ;
        RECT 911.3000 674.8350 913.3000 676.8350 ;
        RECT 935.7500 667.7400 937.7500 669.7400 ;
        RECT 927.6000 667.7400 929.6000 669.7400 ;
        RECT 919.4500 667.7400 921.4500 669.7400 ;
        RECT 911.3000 667.7400 913.3000 669.7400 ;
        RECT 911.3000 689.0250 913.3000 691.0250 ;
        RECT 919.4500 689.0250 921.4500 691.0250 ;
        RECT 927.6000 689.0250 929.6000 691.0250 ;
        RECT 935.7500 689.0250 937.7500 691.0250 ;
        RECT 911.3000 696.1200 913.3000 698.1200 ;
        RECT 919.4500 696.1200 921.4500 698.1200 ;
        RECT 927.6000 696.1200 929.6000 698.1200 ;
        RECT 935.7500 696.1200 937.7500 698.1200 ;
        RECT 952.0500 681.9300 954.0500 683.9300 ;
        RECT 960.2000 681.9300 962.2000 683.9300 ;
        RECT 968.3500 681.9300 970.3500 683.9300 ;
        RECT 976.5000 681.9300 978.5000 683.9300 ;
        RECT 976.5000 674.8350 978.5000 676.8350 ;
        RECT 968.3500 674.8350 970.3500 676.8350 ;
        RECT 960.2000 674.8350 962.2000 676.8350 ;
        RECT 952.0500 674.8350 954.0500 676.8350 ;
        RECT 976.5000 667.7400 978.5000 669.7400 ;
        RECT 968.3500 667.7400 970.3500 669.7400 ;
        RECT 960.2000 667.7400 962.2000 669.7400 ;
        RECT 952.0500 667.7400 954.0500 669.7400 ;
        RECT 952.0500 689.0250 954.0500 691.0250 ;
        RECT 960.2000 689.0250 962.2000 691.0250 ;
        RECT 968.3500 689.0250 970.3500 691.0250 ;
        RECT 976.5000 689.0250 978.5000 691.0250 ;
        RECT 952.0500 696.1200 954.0500 698.1200 ;
        RECT 960.2000 696.1200 962.2000 698.1200 ;
        RECT 968.3500 696.1200 970.3500 698.1200 ;
        RECT 976.5000 696.1200 978.5000 698.1200 ;
        RECT 1049.8500 561.3150 1051.8500 563.3150 ;
        RECT 1049.8500 568.4100 1051.8500 570.4100 ;
        RECT 1049.8500 575.5050 1051.8500 577.5050 ;
        RECT 1049.8500 582.6000 1051.8500 584.6000 ;
        RECT 1049.8500 589.6950 1051.8500 591.6950 ;
        RECT 1049.8500 596.7900 1051.8500 598.7900 ;
        RECT 1049.8500 603.8850 1051.8500 605.8850 ;
        RECT 1049.8500 610.9800 1051.8500 612.9800 ;
        RECT 1049.8500 618.0750 1051.8500 620.0750 ;
        RECT 1049.8500 625.1700 1051.8500 627.1700 ;
        RECT 984.6500 575.5050 986.6500 577.5050 ;
        RECT 992.8000 575.5050 994.8000 577.5050 ;
        RECT 1000.9500 575.5050 1002.9500 577.5050 ;
        RECT 1009.1000 575.5050 1011.1000 577.5050 ;
        RECT 1009.1000 568.4100 1011.1000 570.4100 ;
        RECT 1000.9500 568.4100 1002.9500 570.4100 ;
        RECT 992.8000 568.4100 994.8000 570.4100 ;
        RECT 984.6500 568.4100 986.6500 570.4100 ;
        RECT 1009.1000 561.3150 1011.1000 563.3150 ;
        RECT 1000.9500 561.3150 1002.9500 563.3150 ;
        RECT 992.8000 561.3150 994.8000 563.3150 ;
        RECT 984.6500 561.3150 986.6500 563.3150 ;
        RECT 984.6500 582.6000 986.6500 584.6000 ;
        RECT 992.8000 582.6000 994.8000 584.6000 ;
        RECT 1000.9500 582.6000 1002.9500 584.6000 ;
        RECT 1009.1000 582.6000 1011.1000 584.6000 ;
        RECT 984.6500 589.6950 986.6500 591.6950 ;
        RECT 992.8000 589.6950 994.8000 591.6950 ;
        RECT 1000.9500 589.6950 1002.9500 591.6950 ;
        RECT 1009.1000 589.6950 1011.1000 591.6950 ;
        RECT 1017.2500 575.5050 1019.2500 577.5050 ;
        RECT 1025.4000 575.5050 1027.4000 577.5050 ;
        RECT 1033.5500 575.5050 1035.5500 577.5050 ;
        RECT 1041.7000 575.5050 1043.7000 577.5050 ;
        RECT 1041.7000 568.4100 1043.7000 570.4100 ;
        RECT 1033.5500 568.4100 1035.5500 570.4100 ;
        RECT 1025.4000 568.4100 1027.4000 570.4100 ;
        RECT 1017.2500 568.4100 1019.2500 570.4100 ;
        RECT 1041.7000 561.3150 1043.7000 563.3150 ;
        RECT 1033.5500 561.3150 1035.5500 563.3150 ;
        RECT 1025.4000 561.3150 1027.4000 563.3150 ;
        RECT 1017.2500 561.3150 1019.2500 563.3150 ;
        RECT 1017.2500 582.6000 1019.2500 584.6000 ;
        RECT 1025.4000 582.6000 1027.4000 584.6000 ;
        RECT 1033.5500 582.6000 1035.5500 584.6000 ;
        RECT 1041.7000 582.6000 1043.7000 584.6000 ;
        RECT 1017.2500 589.6950 1019.2500 591.6950 ;
        RECT 1025.4000 589.6950 1027.4000 591.6950 ;
        RECT 1033.5500 589.6950 1035.5500 591.6950 ;
        RECT 1041.7000 589.6950 1043.7000 591.6950 ;
        RECT 984.6500 610.9800 986.6500 612.9800 ;
        RECT 992.8000 610.9800 994.8000 612.9800 ;
        RECT 1000.9500 610.9800 1002.9500 612.9800 ;
        RECT 1009.1000 610.9800 1011.1000 612.9800 ;
        RECT 1009.1000 603.8850 1011.1000 605.8850 ;
        RECT 1000.9500 603.8850 1002.9500 605.8850 ;
        RECT 992.8000 603.8850 994.8000 605.8850 ;
        RECT 984.6500 603.8850 986.6500 605.8850 ;
        RECT 1009.1000 596.7900 1011.1000 598.7900 ;
        RECT 1000.9500 596.7900 1002.9500 598.7900 ;
        RECT 992.8000 596.7900 994.8000 598.7900 ;
        RECT 984.6500 596.7900 986.6500 598.7900 ;
        RECT 984.6500 618.0750 986.6500 620.0750 ;
        RECT 992.8000 618.0750 994.8000 620.0750 ;
        RECT 1000.9500 618.0750 1002.9500 620.0750 ;
        RECT 1009.1000 618.0750 1011.1000 620.0750 ;
        RECT 984.6500 625.1700 986.6500 627.1700 ;
        RECT 992.8000 625.1700 994.8000 627.1700 ;
        RECT 1000.9500 625.1700 1002.9500 627.1700 ;
        RECT 1009.1000 625.1700 1011.1000 627.1700 ;
        RECT 1017.2500 610.9800 1019.2500 612.9800 ;
        RECT 1025.4000 610.9800 1027.4000 612.9800 ;
        RECT 1033.5500 610.9800 1035.5500 612.9800 ;
        RECT 1041.7000 610.9800 1043.7000 612.9800 ;
        RECT 1041.7000 603.8850 1043.7000 605.8850 ;
        RECT 1033.5500 603.8850 1035.5500 605.8850 ;
        RECT 1025.4000 603.8850 1027.4000 605.8850 ;
        RECT 1017.2500 603.8850 1019.2500 605.8850 ;
        RECT 1041.7000 596.7900 1043.7000 598.7900 ;
        RECT 1033.5500 596.7900 1035.5500 598.7900 ;
        RECT 1025.4000 596.7900 1027.4000 598.7900 ;
        RECT 1017.2500 596.7900 1019.2500 598.7900 ;
        RECT 1017.2500 618.0750 1019.2500 620.0750 ;
        RECT 1025.4000 618.0750 1027.4000 620.0750 ;
        RECT 1033.5500 618.0750 1035.5500 620.0750 ;
        RECT 1041.7000 618.0750 1043.7000 620.0750 ;
        RECT 1017.2500 625.1700 1019.2500 627.1700 ;
        RECT 1025.4000 625.1700 1027.4000 627.1700 ;
        RECT 1033.5500 625.1700 1035.5500 627.1700 ;
        RECT 1041.7000 625.1700 1043.7000 627.1700 ;
        RECT 1074.0000 575.5050 1076.0000 577.5050 ;
        RECT 1058.0000 575.5050 1060.0000 577.5050 ;
        RECT 1058.0000 568.4100 1060.0000 570.4100 ;
        RECT 1058.0000 561.3150 1060.0000 563.3150 ;
        RECT 1074.0000 568.4100 1076.0000 570.4100 ;
        RECT 1074.0000 561.3150 1076.0000 563.3150 ;
        RECT 1058.0000 589.6950 1060.0000 591.6950 ;
        RECT 1058.0000 582.6000 1060.0000 584.6000 ;
        RECT 1074.0000 582.6000 1076.0000 584.6000 ;
        RECT 1074.0000 589.6950 1076.0000 591.6950 ;
        RECT 1112.0000 575.5050 1114.0000 577.5050 ;
        RECT 1112.0000 568.4100 1114.0000 570.4100 ;
        RECT 1112.0000 561.3150 1114.0000 563.3150 ;
        RECT 1112.0000 582.6000 1114.0000 584.6000 ;
        RECT 1112.0000 589.6950 1114.0000 591.6950 ;
        RECT 1074.0000 610.9800 1076.0000 612.9800 ;
        RECT 1058.0000 610.9800 1060.0000 612.9800 ;
        RECT 1058.0000 603.8850 1060.0000 605.8850 ;
        RECT 1058.0000 596.7900 1060.0000 598.7900 ;
        RECT 1074.0000 603.8850 1076.0000 605.8850 ;
        RECT 1074.0000 596.7900 1076.0000 598.7900 ;
        RECT 1058.0000 618.0750 1060.0000 620.0750 ;
        RECT 1058.0000 625.1700 1060.0000 627.1700 ;
        RECT 1074.0000 618.0750 1076.0000 620.0750 ;
        RECT 1074.0000 625.1700 1076.0000 627.1700 ;
        RECT 1112.0000 610.9800 1114.0000 612.9800 ;
        RECT 1112.0000 596.7900 1114.0000 598.7900 ;
        RECT 1112.0000 603.8850 1114.0000 605.8850 ;
        RECT 1112.0000 618.0750 1114.0000 620.0750 ;
        RECT 1112.0000 625.1700 1114.0000 627.1700 ;
        RECT 1049.8500 632.2650 1051.8500 634.2650 ;
        RECT 1049.8500 639.3600 1051.8500 641.3600 ;
        RECT 1049.8500 646.4550 1051.8500 648.4550 ;
        RECT 1049.8500 653.5500 1051.8500 655.5500 ;
        RECT 1049.8500 660.6450 1051.8500 662.6450 ;
        RECT 1049.8500 667.7400 1051.8500 669.7400 ;
        RECT 1049.8500 674.8350 1051.8500 676.8350 ;
        RECT 1049.8500 681.9300 1051.8500 683.9300 ;
        RECT 1049.8500 689.0250 1051.8500 691.0250 ;
        RECT 1049.8500 696.1200 1051.8500 698.1200 ;
        RECT 984.6500 646.4550 986.6500 648.4550 ;
        RECT 992.8000 646.4550 994.8000 648.4550 ;
        RECT 1000.9500 646.4550 1002.9500 648.4550 ;
        RECT 1009.1000 646.4550 1011.1000 648.4550 ;
        RECT 1009.1000 639.3600 1011.1000 641.3600 ;
        RECT 1000.9500 639.3600 1002.9500 641.3600 ;
        RECT 992.8000 639.3600 994.8000 641.3600 ;
        RECT 984.6500 639.3600 986.6500 641.3600 ;
        RECT 1009.1000 632.2650 1011.1000 634.2650 ;
        RECT 1000.9500 632.2650 1002.9500 634.2650 ;
        RECT 992.8000 632.2650 994.8000 634.2650 ;
        RECT 984.6500 632.2650 986.6500 634.2650 ;
        RECT 984.6500 653.5500 986.6500 655.5500 ;
        RECT 992.8000 653.5500 994.8000 655.5500 ;
        RECT 1000.9500 653.5500 1002.9500 655.5500 ;
        RECT 1009.1000 653.5500 1011.1000 655.5500 ;
        RECT 984.6500 660.6450 986.6500 662.6450 ;
        RECT 992.8000 660.6450 994.8000 662.6450 ;
        RECT 1000.9500 660.6450 1002.9500 662.6450 ;
        RECT 1009.1000 660.6450 1011.1000 662.6450 ;
        RECT 1017.2500 646.4550 1019.2500 648.4550 ;
        RECT 1025.4000 646.4550 1027.4000 648.4550 ;
        RECT 1033.5500 646.4550 1035.5500 648.4550 ;
        RECT 1041.7000 646.4550 1043.7000 648.4550 ;
        RECT 1041.7000 639.3600 1043.7000 641.3600 ;
        RECT 1033.5500 639.3600 1035.5500 641.3600 ;
        RECT 1025.4000 639.3600 1027.4000 641.3600 ;
        RECT 1017.2500 639.3600 1019.2500 641.3600 ;
        RECT 1041.7000 632.2650 1043.7000 634.2650 ;
        RECT 1033.5500 632.2650 1035.5500 634.2650 ;
        RECT 1025.4000 632.2650 1027.4000 634.2650 ;
        RECT 1017.2500 632.2650 1019.2500 634.2650 ;
        RECT 1017.2500 653.5500 1019.2500 655.5500 ;
        RECT 1025.4000 653.5500 1027.4000 655.5500 ;
        RECT 1033.5500 653.5500 1035.5500 655.5500 ;
        RECT 1041.7000 653.5500 1043.7000 655.5500 ;
        RECT 1017.2500 660.6450 1019.2500 662.6450 ;
        RECT 1025.4000 660.6450 1027.4000 662.6450 ;
        RECT 1033.5500 660.6450 1035.5500 662.6450 ;
        RECT 1041.7000 660.6450 1043.7000 662.6450 ;
        RECT 984.6500 681.9300 986.6500 683.9300 ;
        RECT 992.8000 681.9300 994.8000 683.9300 ;
        RECT 1000.9500 681.9300 1002.9500 683.9300 ;
        RECT 1009.1000 681.9300 1011.1000 683.9300 ;
        RECT 1009.1000 674.8350 1011.1000 676.8350 ;
        RECT 1000.9500 674.8350 1002.9500 676.8350 ;
        RECT 992.8000 674.8350 994.8000 676.8350 ;
        RECT 984.6500 674.8350 986.6500 676.8350 ;
        RECT 1009.1000 667.7400 1011.1000 669.7400 ;
        RECT 1000.9500 667.7400 1002.9500 669.7400 ;
        RECT 992.8000 667.7400 994.8000 669.7400 ;
        RECT 984.6500 667.7400 986.6500 669.7400 ;
        RECT 984.6500 689.0250 986.6500 691.0250 ;
        RECT 992.8000 689.0250 994.8000 691.0250 ;
        RECT 1000.9500 689.0250 1002.9500 691.0250 ;
        RECT 1009.1000 689.0250 1011.1000 691.0250 ;
        RECT 984.6500 696.1200 986.6500 698.1200 ;
        RECT 992.8000 696.1200 994.8000 698.1200 ;
        RECT 1000.9500 696.1200 1002.9500 698.1200 ;
        RECT 1009.1000 696.1200 1011.1000 698.1200 ;
        RECT 1017.2500 681.9300 1019.2500 683.9300 ;
        RECT 1025.4000 681.9300 1027.4000 683.9300 ;
        RECT 1033.5500 681.9300 1035.5500 683.9300 ;
        RECT 1041.7000 681.9300 1043.7000 683.9300 ;
        RECT 1041.7000 674.8350 1043.7000 676.8350 ;
        RECT 1033.5500 674.8350 1035.5500 676.8350 ;
        RECT 1025.4000 674.8350 1027.4000 676.8350 ;
        RECT 1017.2500 674.8350 1019.2500 676.8350 ;
        RECT 1041.7000 667.7400 1043.7000 669.7400 ;
        RECT 1033.5500 667.7400 1035.5500 669.7400 ;
        RECT 1025.4000 667.7400 1027.4000 669.7400 ;
        RECT 1017.2500 667.7400 1019.2500 669.7400 ;
        RECT 1017.2500 689.0250 1019.2500 691.0250 ;
        RECT 1025.4000 689.0250 1027.4000 691.0250 ;
        RECT 1033.5500 689.0250 1035.5500 691.0250 ;
        RECT 1041.7000 689.0250 1043.7000 691.0250 ;
        RECT 1017.2500 696.1200 1019.2500 698.1200 ;
        RECT 1025.4000 696.1200 1027.4000 698.1200 ;
        RECT 1033.5500 696.1200 1035.5500 698.1200 ;
        RECT 1041.7000 696.1200 1043.7000 698.1200 ;
        RECT 1074.0000 646.4550 1076.0000 648.4550 ;
        RECT 1058.0000 646.4550 1060.0000 648.4550 ;
        RECT 1058.0000 639.3600 1060.0000 641.3600 ;
        RECT 1058.0000 632.2650 1060.0000 634.2650 ;
        RECT 1074.0000 632.2650 1076.0000 634.2650 ;
        RECT 1074.0000 639.3600 1076.0000 641.3600 ;
        RECT 1058.0000 660.6450 1060.0000 662.6450 ;
        RECT 1058.0000 653.5500 1060.0000 655.5500 ;
        RECT 1074.0000 660.6450 1076.0000 662.6450 ;
        RECT 1074.0000 653.5500 1076.0000 655.5500 ;
        RECT 1112.0000 646.4550 1114.0000 648.4550 ;
        RECT 1112.0000 632.2650 1114.0000 634.2650 ;
        RECT 1112.0000 639.3600 1114.0000 641.3600 ;
        RECT 1112.0000 653.5500 1114.0000 655.5500 ;
        RECT 1112.0000 660.6450 1114.0000 662.6450 ;
        RECT 1074.0000 681.9300 1076.0000 683.9300 ;
        RECT 1058.0000 681.9300 1060.0000 683.9300 ;
        RECT 1058.0000 674.8350 1060.0000 676.8350 ;
        RECT 1058.0000 667.7400 1060.0000 669.7400 ;
        RECT 1074.0000 667.7400 1076.0000 669.7400 ;
        RECT 1074.0000 674.8350 1076.0000 676.8350 ;
        RECT 1058.0000 696.1200 1060.0000 698.1200 ;
        RECT 1058.0000 689.0250 1060.0000 691.0250 ;
        RECT 1074.0000 689.0250 1076.0000 691.0250 ;
        RECT 1074.0000 696.1200 1076.0000 698.1200 ;
        RECT 1112.0000 681.9300 1114.0000 683.9300 ;
        RECT 1112.0000 667.7400 1114.0000 669.7400 ;
        RECT 1112.0000 674.8350 1114.0000 676.8350 ;
        RECT 1112.0000 689.0250 1114.0000 691.0250 ;
        RECT 1112.0000 696.1200 1114.0000 698.1200 ;
        RECT 846.1000 703.2150 848.1000 705.2150 ;
        RECT 854.2500 703.2150 856.2500 705.2150 ;
        RECT 862.4000 703.2150 864.4000 705.2150 ;
        RECT 870.5500 703.2150 872.5500 705.2150 ;
        RECT 878.7000 703.2150 880.7000 705.2150 ;
        RECT 886.8500 703.2150 888.8500 705.2150 ;
        RECT 895.0000 703.2150 897.0000 705.2150 ;
        RECT 903.1500 703.2150 905.1500 705.2150 ;
        RECT 952.0500 703.2150 954.0500 705.2150 ;
        RECT 911.3000 703.2150 913.3000 705.2150 ;
        RECT 919.4500 703.2150 921.4500 705.2150 ;
        RECT 927.6000 703.2150 929.6000 705.2150 ;
        RECT 935.7500 703.2150 937.7500 705.2150 ;
        RECT 943.9000 703.2150 945.9000 705.2150 ;
        RECT 960.2000 703.2150 962.2000 705.2150 ;
        RECT 968.3500 703.2150 970.3500 705.2150 ;
        RECT 976.5000 703.2150 978.5000 705.2150 ;
        RECT 1049.8500 703.2150 1051.8500 705.2150 ;
        RECT 984.6500 703.2150 986.6500 705.2150 ;
        RECT 992.8000 703.2150 994.8000 705.2150 ;
        RECT 1000.9500 703.2150 1002.9500 705.2150 ;
        RECT 1009.1000 703.2150 1011.1000 705.2150 ;
        RECT 1017.2500 703.2150 1019.2500 705.2150 ;
        RECT 1025.4000 703.2150 1027.4000 705.2150 ;
        RECT 1033.5500 703.2150 1035.5500 705.2150 ;
        RECT 1041.7000 703.2150 1043.7000 705.2150 ;
        RECT 1074.0000 717.4050 1076.0000 719.4050 ;
        RECT 1058.0000 708.0000 1060.0000 710.0000 ;
        RECT 1058.0000 703.2150 1060.0000 705.2150 ;
        RECT 1074.0000 710.3100 1076.0000 712.3100 ;
        RECT 1074.0000 703.2150 1076.0000 705.2150 ;
        RECT 1074.0000 724.5000 1076.0000 726.0000 ;
        RECT 1112.0000 717.4050 1114.0000 719.4050 ;
        RECT 1112.0000 703.2150 1114.0000 705.2150 ;
        RECT 1112.0000 710.3100 1114.0000 712.3100 ;
        RECT 1112.0000 724.5000 1114.0000 726.5000 ;
        RECT 1112.0000 731.5950 1114.0000 733.5950 ;
        RECT 1112.0000 738.6900 1114.0000 740.6900 ;
        RECT 1112.0000 745.7850 1114.0000 747.7850 ;
        RECT 1112.0000 759.9750 1114.0000 761.9750 ;
        RECT 1112.0000 752.8800 1114.0000 754.8800 ;
        RECT 1112.0000 767.0700 1114.0000 769.0700 ;
        RECT 1112.0000 774.1650 1114.0000 776.1650 ;
        RECT 1112.0000 781.2600 1114.0000 783.2600 ;
        RECT 1112.0000 795.4500 1114.0000 797.4500 ;
        RECT 1112.0000 788.3550 1114.0000 790.3550 ;
        RECT 1112.0000 802.5450 1114.0000 804.5450 ;
        RECT 1112.0000 809.6400 1114.0000 811.6400 ;
        RECT 1112.0000 816.7350 1114.0000 818.7350 ;
        RECT 1112.0000 830.9250 1114.0000 832.9250 ;
        RECT 1112.0000 823.8300 1114.0000 825.8300 ;
        RECT 1112.0000 979.9200 1114.0000 981.9200 ;
        RECT 1112.0000 908.9700 1114.0000 910.9700 ;
        RECT 1112.0000 873.4950 1114.0000 875.4950 ;
        RECT 1112.0000 845.1150 1114.0000 847.1150 ;
        RECT 1112.0000 852.2100 1114.0000 854.2100 ;
        RECT 1112.0000 859.3050 1114.0000 861.3050 ;
        RECT 1112.0000 866.4000 1114.0000 868.4000 ;
        RECT 1112.0000 880.5900 1114.0000 882.5900 ;
        RECT 1112.0000 887.6850 1114.0000 889.6850 ;
        RECT 1112.0000 894.7800 1114.0000 896.7800 ;
        RECT 1112.0000 901.8750 1114.0000 903.8750 ;
        RECT 1112.0000 944.4450 1114.0000 946.4450 ;
        RECT 1112.0000 916.0650 1114.0000 918.0650 ;
        RECT 1112.0000 923.1600 1114.0000 925.1600 ;
        RECT 1112.0000 930.2550 1114.0000 932.2550 ;
        RECT 1112.0000 937.3500 1114.0000 939.3500 ;
        RECT 1112.0000 951.5400 1114.0000 953.5400 ;
        RECT 1112.0000 958.6350 1114.0000 960.6350 ;
        RECT 1112.0000 965.7300 1114.0000 967.7300 ;
        RECT 1112.0000 972.8250 1114.0000 974.8250 ;
        RECT 1112.0000 987.0150 1114.0000 989.0150 ;
        RECT 1112.0000 994.1100 1114.0000 996.1100 ;
        RECT 1112.0000 1001.2050 1114.0000 1003.2050 ;
        RECT 1112.0000 1008.3000 1114.0000 1010.3000 ;
        RECT 1112.0000 1022.4900 1114.0000 1024.4900 ;
        RECT 1112.0000 1015.3950 1114.0000 1017.3950 ;
        RECT 1112.0000 1029.5850 1114.0000 1031.5850 ;
        RECT 1112.0000 1036.6800 1114.0000 1038.6800 ;
        RECT 1112.0000 1043.7750 1114.0000 1045.7750 ;
        RECT 1112.0000 1057.9650 1114.0000 1059.9650 ;
        RECT 1112.0000 1050.8700 1114.0000 1052.8700 ;
        RECT 1112.0000 1065.0600 1114.0000 1067.0600 ;
        RECT 1112.0000 1072.1550 1114.0000 1074.1550 ;
        RECT 1112.0000 1079.2500 1114.0000 1081.2500 ;
        RECT 1112.0000 1100.5350 1114.0000 1102.5350 ;
        RECT 1112.0000 1093.4400 1114.0000 1095.4400 ;
        RECT 1112.0000 1086.3450 1114.0000 1088.3450 ;
        RECT 1112.0000 1107.6300 1114.0000 1109.6300 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'sram_w16_64b'
    PORT
      LAYER M4 ;
        RECT 323.9650 60.0000 325.9650 330.0000 ;
        RECT 306.9350 60.0000 308.9350 330.0000 ;
        RECT 315.4500 60.0000 317.4500 330.0000 ;
        RECT 298.4200 60.0000 300.4200 330.0000 ;
        RECT 289.9050 60.0000 291.9050 330.0000 ;
        RECT 281.3900 60.0000 283.3900 330.0000 ;
        RECT 272.8750 60.0000 274.8750 330.0000 ;
        RECT 264.3600 60.0000 266.3600 330.0000 ;
        RECT 255.8450 60.0000 257.8450 330.0000 ;
        RECT 247.3300 60.0000 249.3300 330.0000 ;
        RECT 238.8150 60.0000 240.8150 330.0000 ;
        RECT 221.7850 60.0000 223.7850 330.0000 ;
        RECT 213.2700 60.0000 215.2700 330.0000 ;
        RECT 204.7550 60.0000 206.7550 330.0000 ;
        RECT 196.2400 60.0000 198.2400 330.0000 ;
        RECT 230.3000 60.0000 232.3000 330.0000 ;
        RECT 187.7250 60.0000 189.7250 330.0000 ;
        RECT 179.2100 60.0000 181.2100 330.0000 ;
        RECT 170.6950 60.0000 172.6950 330.0000 ;
        RECT 162.1800 60.0000 164.1800 330.0000 ;
        RECT 153.6650 60.0000 155.6650 330.0000 ;
        RECT 145.1500 60.0000 147.1500 330.0000 ;
        RECT 136.6350 60.0000 138.6350 330.0000 ;
        RECT 128.1200 60.0000 130.1200 330.0000 ;
        RECT 119.6050 60.0000 121.6050 330.0000 ;
        RECT 111.0900 60.0000 113.0900 330.0000 ;
        RECT 94.0600 60.0000 96.0600 330.0000 ;
        RECT 102.5750 60.0000 104.5750 330.0000 ;
        RECT 60.0000 60.0000 62.0000 330.0000 ;
        RECT 68.5150 60.0000 70.5150 330.0000 ;
        RECT 77.0300 60.0000 79.0300 330.0000 ;
        RECT 85.5450 60.0000 87.5450 330.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16_64b'


# P/G pin shape extracted from block 'sram_w16_64b'
    PORT
      LAYER M4 ;
        RECT 323.9650 410.0000 325.9650 680.0000 ;
        RECT 306.9350 410.0000 308.9350 680.0000 ;
        RECT 315.4500 410.0000 317.4500 680.0000 ;
        RECT 298.4200 410.0000 300.4200 680.0000 ;
        RECT 289.9050 410.0000 291.9050 680.0000 ;
        RECT 281.3900 410.0000 283.3900 680.0000 ;
        RECT 272.8750 410.0000 274.8750 680.0000 ;
        RECT 264.3600 410.0000 266.3600 680.0000 ;
        RECT 255.8450 410.0000 257.8450 680.0000 ;
        RECT 247.3300 410.0000 249.3300 680.0000 ;
        RECT 238.8150 410.0000 240.8150 680.0000 ;
        RECT 221.7850 410.0000 223.7850 680.0000 ;
        RECT 213.2700 410.0000 215.2700 680.0000 ;
        RECT 204.7550 410.0000 206.7550 680.0000 ;
        RECT 196.2400 410.0000 198.2400 680.0000 ;
        RECT 230.3000 410.0000 232.3000 680.0000 ;
        RECT 187.7250 410.0000 189.7250 680.0000 ;
        RECT 179.2100 410.0000 181.2100 680.0000 ;
        RECT 170.6950 410.0000 172.6950 680.0000 ;
        RECT 162.1800 410.0000 164.1800 680.0000 ;
        RECT 153.6650 410.0000 155.6650 680.0000 ;
        RECT 145.1500 410.0000 147.1500 680.0000 ;
        RECT 136.6350 410.0000 138.6350 680.0000 ;
        RECT 128.1200 410.0000 130.1200 680.0000 ;
        RECT 119.6050 410.0000 121.6050 680.0000 ;
        RECT 111.0900 410.0000 113.0900 680.0000 ;
        RECT 94.0600 410.0000 96.0600 680.0000 ;
        RECT 102.5750 410.0000 104.5750 680.0000 ;
        RECT 60.0000 410.0000 62.0000 680.0000 ;
        RECT 68.5150 410.0000 70.5150 680.0000 ;
        RECT 77.0300 410.0000 79.0300 680.0000 ;
        RECT 85.5450 410.0000 87.5450 680.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16_64b'


# P/G pin shape extracted from block 'sram_w16_160b'
    PORT
      LAYER M4 ;
        RECT 479.3500 60.0000 481.3500 710.0000 ;
        RECT 471.2000 60.0000 473.2000 710.0000 ;
        RECT 463.0500 60.0000 465.0500 710.0000 ;
        RECT 454.9000 60.0000 456.9000 710.0000 ;
        RECT 446.7500 60.0000 448.7500 710.0000 ;
        RECT 438.6000 60.0000 440.6000 710.0000 ;
        RECT 430.4500 60.0000 432.4500 710.0000 ;
        RECT 422.3000 60.0000 424.3000 710.0000 ;
        RECT 414.1500 60.0000 416.1500 710.0000 ;
        RECT 495.6500 60.0000 497.6500 710.0000 ;
        RECT 503.8000 60.0000 505.8000 710.0000 ;
        RECT 511.9500 60.0000 513.9500 710.0000 ;
        RECT 520.1000 60.0000 522.1000 710.0000 ;
        RECT 528.2500 60.0000 530.2500 710.0000 ;
        RECT 536.4000 60.0000 538.4000 710.0000 ;
        RECT 544.5500 60.0000 546.5500 710.0000 ;
        RECT 552.7000 60.0000 554.7000 710.0000 ;
        RECT 560.8500 60.0000 562.8500 710.0000 ;
        RECT 487.5000 60.0000 489.5000 710.0000 ;
        RECT 569.0000 60.0000 571.0000 710.0000 ;
        RECT 577.1500 60.0000 579.1500 710.0000 ;
        RECT 585.3000 60.0000 587.3000 710.0000 ;
        RECT 593.4500 60.0000 595.4500 710.0000 ;
        RECT 601.6000 60.0000 603.6000 710.0000 ;
        RECT 609.7500 60.0000 611.7500 710.0000 ;
        RECT 617.9000 60.0000 619.9000 710.0000 ;
        RECT 626.0500 60.0000 628.0500 710.0000 ;
        RECT 634.2000 60.0000 636.2000 710.0000 ;
        RECT 642.3500 60.0000 644.3500 710.0000 ;
        RECT 658.6500 60.0000 660.6500 710.0000 ;
        RECT 666.8000 60.0000 668.8000 710.0000 ;
        RECT 674.9500 60.0000 676.9500 710.0000 ;
        RECT 683.1000 60.0000 685.1000 710.0000 ;
        RECT 691.2500 60.0000 693.2500 710.0000 ;
        RECT 699.4000 60.0000 701.4000 710.0000 ;
        RECT 707.5500 60.0000 709.5500 710.0000 ;
        RECT 715.7000 60.0000 717.7000 710.0000 ;
        RECT 723.8500 60.0000 725.8500 710.0000 ;
        RECT 732.0000 60.0000 734.0000 710.0000 ;
        RECT 650.5000 60.0000 652.5000 710.0000 ;
        RECT 805.3500 60.0000 807.3500 710.0000 ;
        RECT 813.5000 60.0000 815.5000 710.0000 ;
        RECT 797.2000 60.0000 799.2000 710.0000 ;
        RECT 789.0500 60.0000 791.0500 710.0000 ;
        RECT 780.9000 60.0000 782.9000 710.0000 ;
        RECT 772.7500 60.0000 774.7500 710.0000 ;
        RECT 764.6000 60.0000 766.6000 710.0000 ;
        RECT 756.4500 60.0000 758.4500 710.0000 ;
        RECT 748.3000 60.0000 750.3000 710.0000 ;
        RECT 740.1500 60.0000 742.1500 710.0000 ;
        RECT 895.0000 60.0000 897.0000 710.0000 ;
        RECT 886.8500 60.0000 888.8500 710.0000 ;
        RECT 878.7000 60.0000 880.7000 710.0000 ;
        RECT 870.5500 60.0000 872.5500 710.0000 ;
        RECT 862.4000 60.0000 864.4000 710.0000 ;
        RECT 854.2500 60.0000 856.2500 710.0000 ;
        RECT 846.1000 60.0000 848.1000 710.0000 ;
        RECT 837.9500 60.0000 839.9500 710.0000 ;
        RECT 829.8000 60.0000 831.8000 710.0000 ;
        RECT 821.6500 60.0000 823.6500 710.0000 ;
        RECT 976.5000 60.0000 978.5000 710.0000 ;
        RECT 968.3500 60.0000 970.3500 710.0000 ;
        RECT 960.2000 60.0000 962.2000 710.0000 ;
        RECT 952.0500 60.0000 954.0500 710.0000 ;
        RECT 943.9000 60.0000 945.9000 710.0000 ;
        RECT 935.7500 60.0000 937.7500 710.0000 ;
        RECT 927.6000 60.0000 929.6000 710.0000 ;
        RECT 919.4500 60.0000 921.4500 710.0000 ;
        RECT 911.3000 60.0000 913.3000 710.0000 ;
        RECT 903.1500 60.0000 905.1500 710.0000 ;
        RECT 1058.0000 60.0000 1060.0000 710.0000 ;
        RECT 1049.8500 60.0000 1051.8500 710.0000 ;
        RECT 1041.7000 60.0000 1043.7000 710.0000 ;
        RECT 1033.5500 60.0000 1035.5500 710.0000 ;
        RECT 1025.4000 60.0000 1027.4000 710.0000 ;
        RECT 1017.2500 60.0000 1019.2500 710.0000 ;
        RECT 1009.1000 60.0000 1011.1000 710.0000 ;
        RECT 1000.9500 60.0000 1002.9500 710.0000 ;
        RECT 992.8000 60.0000 994.8000 710.0000 ;
        RECT 984.6500 60.0000 986.6500 710.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16_160b'

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 1114.1000 279.6100 1116.1000 281.6100 ;
        RECT 1114.5000 2.0000 1116.5000 39.3800 ;
        RECT 1114.5000 17.0950 1116.5000 19.0950 ;
        RECT 1114.5000 2.0000 1116.5000 18.0950 ;
        RECT 1114.5000 2.0000 1116.5000 32.2850 ;
        RECT 1114.5000 2.0000 1116.5000 25.1900 ;
        RECT 1114.5000 24.1900 1116.5000 26.1900 ;
        RECT 1114.5000 31.2850 1116.5000 33.2850 ;
        RECT 1114.5000 38.3800 1116.5000 40.3800 ;
        RECT 1114.1000 46.4750 1116.1000 48.0000 ;
        RECT 1114.1000 45.4750 1116.1000 47.4750 ;
        RECT 1114.1000 59.6650 1116.1000 61.6650 ;
        RECT 1114.1000 52.5700 1116.1000 54.5700 ;
        RECT 1114.1000 53.5700 1116.1000 54.0000 ;
        RECT 1114.1000 60.6650 1116.1000 61.2000 ;
        RECT 1114.1000 67.7600 1116.1000 68.2000 ;
        RECT 1114.1000 66.7600 1116.1000 68.7600 ;
        RECT 1114.1000 74.8550 1116.1000 75.4000 ;
        RECT 1114.1000 73.8550 1116.1000 75.8550 ;
        RECT 1114.1000 80.9500 1116.1000 82.9500 ;
        RECT 1114.1000 81.9500 1116.1000 82.4000 ;
        RECT 1114.1000 95.1400 1116.1000 97.1400 ;
        RECT 1114.1000 96.1400 1116.1000 96.6000 ;
        RECT 1114.1000 88.0450 1116.1000 90.0450 ;
        RECT 1114.1000 89.0450 1116.1000 89.6000 ;
        RECT 1114.1000 102.2350 1116.1000 104.2350 ;
        RECT 1114.1000 103.2350 1116.1000 103.8000 ;
        RECT 1114.1000 110.3300 1116.1000 110.8000 ;
        RECT 1114.1000 109.3300 1116.1000 111.3300 ;
        RECT 1114.1000 117.4250 1116.1000 118.0000 ;
        RECT 1114.1000 116.4250 1116.1000 118.4250 ;
        RECT 1114.1000 130.6150 1116.1000 132.6150 ;
        RECT 1114.1000 124.5200 1116.1000 125.0000 ;
        RECT 1114.1000 123.5200 1116.1000 125.5200 ;
        RECT 1114.1000 131.6150 1116.1000 132.2000 ;
        RECT 1114.1000 137.7100 1116.1000 139.7100 ;
        RECT 1114.1000 138.7100 1116.1000 139.2000 ;
        RECT 1114.1000 208.6600 1116.1000 210.6600 ;
        RECT 1114.1000 209.6600 1116.1000 210.2000 ;
        RECT 1114.1000 173.1850 1116.1000 175.1850 ;
        RECT 1114.1000 144.8050 1116.1000 146.8050 ;
        RECT 1114.1000 145.8050 1116.1000 146.4000 ;
        RECT 1114.1000 151.9000 1116.1000 153.9000 ;
        RECT 1114.1000 152.9000 1116.1000 153.4000 ;
        RECT 1114.1000 166.0900 1116.1000 168.0900 ;
        RECT 1114.1000 158.9950 1116.1000 160.9950 ;
        RECT 1114.1000 159.9950 1116.1000 160.4000 ;
        RECT 1114.1000 174.1850 1116.1000 174.6000 ;
        RECT 1114.1000 167.0900 1116.1000 167.6000 ;
        RECT 1114.1000 180.2800 1116.1000 182.2800 ;
        RECT 1114.1000 181.2800 1116.1000 181.8000 ;
        RECT 1114.1000 187.3750 1116.1000 189.3750 ;
        RECT 1114.1000 188.3750 1116.1000 188.8000 ;
        RECT 1114.1000 194.4700 1116.1000 196.4700 ;
        RECT 1114.1000 195.4700 1116.1000 196.0000 ;
        RECT 1114.1000 201.5650 1116.1000 203.5650 ;
        RECT 1114.1000 202.5650 1116.1000 203.0000 ;
        RECT 1114.1000 244.1350 1116.1000 246.1350 ;
        RECT 1114.1000 215.7550 1116.1000 217.7550 ;
        RECT 1114.1000 216.7550 1116.1000 217.2000 ;
        RECT 1114.1000 222.8500 1116.1000 224.8500 ;
        RECT 1114.1000 223.8500 1116.1000 224.4000 ;
        RECT 1114.1000 229.9450 1116.1000 231.9450 ;
        RECT 1114.1000 230.9450 1116.1000 231.4000 ;
        RECT 1114.1000 237.0400 1116.1000 239.0400 ;
        RECT 1114.1000 238.0400 1116.1000 238.6000 ;
        RECT 1114.1000 251.2300 1116.1000 253.2300 ;
        RECT 1114.1000 252.2300 1116.1000 252.8000 ;
        RECT 1114.1000 245.1350 1116.1000 245.6000 ;
        RECT 1114.1000 258.3250 1116.1000 260.3250 ;
        RECT 1114.1000 259.3250 1116.1000 259.8000 ;
        RECT 1114.1000 266.4200 1116.1000 267.4000 ;
        RECT 1114.1000 265.4200 1116.1000 267.4200 ;
        RECT 1114.1000 272.5150 1116.1000 274.5150 ;
        RECT 1114.1000 273.5150 1116.1000 274.6000 ;
        RECT 1114.1000 287.7050 1116.1000 288.2000 ;
        RECT 1114.1000 286.7050 1116.1000 288.7050 ;
        RECT 1114.1000 280.6100 1116.1000 281.8000 ;
        RECT 1114.1000 294.8000 1116.1000 295.4000 ;
        RECT 1114.1000 293.8000 1116.1000 295.8000 ;
        RECT 1114.1000 300.8950 1116.1000 302.8950 ;
        RECT 1114.1000 301.8950 1116.1000 302.4000 ;
        RECT 1114.1000 308.9900 1116.1000 309.4000 ;
        RECT 1114.1000 307.9900 1116.1000 309.9900 ;
        RECT 1114.1000 322.1800 1116.1000 324.1800 ;
        RECT 1114.1000 315.0850 1116.1000 317.0850 ;
        RECT 1114.1000 316.0850 1116.1000 316.6000 ;
        RECT 1114.1000 323.1800 1116.1000 323.6000 ;
        RECT 1114.1000 330.2750 1116.1000 330.8000 ;
        RECT 1114.1000 329.2750 1116.1000 331.2750 ;
        RECT 1114.1000 336.3700 1116.1000 338.3700 ;
        RECT 1114.1000 337.3700 1116.1000 337.8000 ;
        RECT 1114.1000 343.4650 1116.1000 345.4650 ;
        RECT 1114.1000 344.4650 1116.1000 345.0000 ;
        RECT 1071.0000 373.8000 1073.0000 375.8000 ;
        RECT 1114.1000 357.6550 1116.1000 359.6550 ;
        RECT 1114.1000 358.6550 1116.1000 359.2000 ;
        RECT 1114.1000 351.5600 1116.1000 352.0000 ;
        RECT 1114.1000 350.5600 1116.1000 352.5600 ;
        RECT 1114.1000 364.7500 1116.1000 366.7500 ;
        RECT 1114.1000 365.7500 1116.1000 366.2000 ;
        RECT 1114.1000 371.8450 1116.1000 373.8450 ;
        RECT 1114.1000 372.8450 1116.1000 374.6000 ;
        RECT 1114.1000 393.1300 1116.1000 395.1300 ;
        RECT 1114.1000 386.0350 1116.1000 388.0350 ;
        RECT 1114.1000 387.0350 1116.1000 387.6000 ;
        RECT 1114.1000 394.1300 1116.1000 394.8000 ;
        RECT 1114.1000 400.2250 1116.1000 402.2250 ;
        RECT 1114.1000 401.2250 1116.1000 401.8000 ;
        RECT 1114.1000 407.3200 1116.1000 409.3200 ;
        RECT 1114.1000 408.3200 1116.1000 408.8000 ;
        RECT 1114.1000 414.4150 1116.1000 416.4150 ;
        RECT 1114.1000 415.4150 1116.1000 416.0000 ;
        RECT 1114.1000 435.7000 1116.1000 437.7000 ;
        RECT 1114.1000 428.6050 1116.1000 430.6050 ;
        RECT 1114.1000 421.5100 1116.1000 423.5100 ;
        RECT 1114.1000 422.5100 1116.1000 423.0000 ;
        RECT 1114.1000 429.6050 1116.1000 430.2000 ;
        RECT 1114.1000 436.7000 1116.1000 437.2000 ;
        RECT 1114.1000 442.7950 1116.1000 444.7950 ;
        RECT 1114.1000 443.7950 1116.1000 444.2000 ;
        RECT 1114.1000 449.8900 1116.1000 451.8900 ;
        RECT 1114.1000 450.8900 1116.1000 451.4000 ;
        RECT 1114.1000 471.1750 1116.1000 473.1750 ;
        RECT 1114.1000 472.1750 1116.1000 472.6000 ;
        RECT 1114.1000 456.9850 1116.1000 458.9850 ;
        RECT 1114.1000 457.9850 1116.1000 458.4000 ;
        RECT 1114.1000 464.0800 1116.1000 466.0800 ;
        RECT 1114.1000 465.0800 1116.1000 465.6000 ;
        RECT 1114.1000 478.2700 1116.1000 480.2700 ;
        RECT 1114.1000 479.2700 1116.1000 479.8000 ;
        RECT 1114.1000 485.3650 1116.1000 487.3650 ;
        RECT 1114.1000 486.3650 1116.1000 486.8000 ;
        RECT 1114.1000 506.6500 1116.1000 508.6500 ;
        RECT 1114.1000 492.4600 1116.1000 494.4600 ;
        RECT 1114.1000 493.4600 1116.1000 494.0000 ;
        RECT 1114.1000 499.5550 1116.1000 501.5550 ;
        RECT 1114.1000 500.5550 1116.1000 501.0000 ;
        RECT 1114.1000 513.7450 1116.1000 515.7450 ;
        RECT 1114.1000 514.7450 1116.1000 515.8000 ;
        RECT 1114.1000 507.6500 1116.1000 508.2000 ;
        RECT 1114.1000 521.8400 1116.1000 523.0000 ;
        RECT 1114.1000 520.8400 1116.1000 522.8400 ;
        RECT 1114.1000 542.1250 1116.1000 544.1250 ;
        RECT 1114.1000 527.9350 1116.1000 529.9350 ;
        RECT 1114.1000 528.9350 1116.1000 529.4000 ;
        RECT 1114.1000 535.0300 1116.1000 537.0300 ;
        RECT 1114.1000 536.0300 1116.1000 536.6000 ;
        RECT 1114.1000 543.1250 1116.1000 543.6000 ;
        RECT 1114.1000 549.2200 1116.1000 551.2200 ;
        RECT 1114.1000 550.2200 1116.1000 550.8000 ;
        RECT 1114.1000 557.3150 1116.1000 557.8000 ;
        RECT 1114.1000 556.3150 1116.1000 558.3150 ;
        RECT 1114.1000 698.2150 1116.1000 700.2150 ;
        RECT 1114.1000 564.4100 1116.1000 565.0000 ;
        RECT 1114.1000 563.4100 1116.1000 565.4100 ;
        RECT 1114.1000 570.5050 1116.1000 572.5050 ;
        RECT 1114.1000 571.5050 1116.1000 572.0000 ;
        RECT 1114.1000 584.6950 1116.1000 586.6950 ;
        RECT 1114.1000 577.6000 1116.1000 579.6000 ;
        RECT 1114.1000 578.6000 1116.1000 579.2000 ;
        RECT 1114.1000 585.6950 1116.1000 586.2000 ;
        RECT 1114.1000 591.7900 1116.1000 593.7900 ;
        RECT 1114.1000 592.7900 1116.1000 593.2000 ;
        RECT 1114.1000 598.8850 1116.1000 600.8850 ;
        RECT 1114.1000 599.8850 1116.1000 600.4000 ;
        RECT 1114.1000 606.9800 1116.1000 607.4000 ;
        RECT 1114.1000 605.9800 1116.1000 607.9800 ;
        RECT 1114.1000 620.1700 1116.1000 622.1700 ;
        RECT 1114.1000 621.1700 1116.1000 621.6000 ;
        RECT 1114.1000 613.0750 1116.1000 615.0750 ;
        RECT 1114.1000 614.0750 1116.1000 614.6000 ;
        RECT 1114.1000 628.2650 1116.1000 628.8000 ;
        RECT 1114.1000 627.2650 1116.1000 629.2650 ;
        RECT 1114.1000 634.3600 1116.1000 636.3600 ;
        RECT 1114.1000 635.3600 1116.1000 635.8000 ;
        RECT 1114.1000 641.4550 1116.1000 643.4550 ;
        RECT 1114.1000 642.4550 1116.1000 643.0000 ;
        RECT 1114.1000 655.6450 1116.1000 657.6450 ;
        RECT 1114.1000 648.5500 1116.1000 650.5500 ;
        RECT 1114.1000 649.5500 1116.1000 650.0000 ;
        RECT 1114.1000 656.6450 1116.1000 657.2000 ;
        RECT 1114.1000 662.7400 1116.1000 664.7400 ;
        RECT 1114.1000 663.7400 1116.1000 664.2000 ;
        RECT 1114.1000 669.8350 1116.1000 671.8350 ;
        RECT 1114.1000 670.8350 1116.1000 671.4000 ;
        RECT 1114.1000 676.9300 1116.1000 678.9300 ;
        RECT 1114.1000 677.9300 1116.1000 678.4000 ;
        RECT 1114.1000 691.1200 1116.1000 693.1200 ;
        RECT 1114.1000 684.0250 1116.1000 686.0250 ;
        RECT 1114.1000 685.0250 1116.1000 685.6000 ;
        RECT 1114.1000 692.1200 1116.1000 692.6000 ;
        RECT 1114.1000 699.2150 1116.1000 699.8000 ;
        RECT 1114.5000 769.1650 1116.5000 771.1650 ;
        RECT 1114.5000 722.0000 1116.5000 784.3550 ;
        RECT 1114.5000 722.0000 1116.5000 777.2600 ;
        RECT 1114.5000 722.0000 1116.5000 770.1650 ;
        RECT 1114.5000 722.0000 1116.5000 763.0700 ;
        RECT 1114.5000 722.0000 1116.5000 755.9750 ;
        RECT 1114.5000 722.0000 1116.5000 748.8800 ;
        RECT 1114.5000 722.0000 1116.5000 741.7850 ;
        RECT 1114.5000 733.6900 1116.5000 735.6900 ;
        RECT 1114.1000 705.3100 1116.1000 707.3100 ;
        RECT 1114.1000 706.3100 1116.1000 706.8000 ;
        RECT 1114.1000 712.4050 1116.1000 714.4050 ;
        RECT 1114.1000 713.4050 1116.1000 714.0000 ;
        RECT 1114.5000 722.0000 1116.5000 734.6900 ;
        RECT 1114.5000 722.0000 1116.5000 727.5950 ;
        RECT 1114.1000 719.5000 1116.1000 721.5000 ;
        RECT 1114.1000 720.5000 1116.1000 721.0000 ;
        RECT 1114.5000 726.5950 1116.5000 728.5950 ;
        RECT 1114.5000 740.7850 1116.5000 742.7850 ;
        RECT 1114.5000 747.8800 1116.5000 749.8800 ;
        RECT 1114.5000 754.9750 1116.5000 756.9750 ;
        RECT 1114.5000 762.0700 1116.5000 764.0700 ;
        RECT 1114.5000 776.2600 1116.5000 778.2600 ;
        RECT 1114.5000 783.3550 1116.5000 785.3550 ;
        RECT 1114.5000 1011.3950 1116.5000 1117.9000 ;
        RECT 1114.5000 1018.4900 1116.5000 1117.9000 ;
        RECT 1114.5000 1025.5850 1116.5000 1117.9000 ;
        RECT 1114.5000 1032.6800 1116.5000 1117.9000 ;
        RECT 1114.5000 1039.7750 1116.5000 1117.9000 ;
        RECT 1114.5000 1046.8700 1116.5000 1117.9000 ;
        RECT 1114.5000 1010.3950 1116.5000 1012.3950 ;
        RECT 1114.5000 1031.6800 1116.5000 1033.6800 ;
        RECT 1114.5000 1017.4900 1116.5000 1019.4900 ;
        RECT 1114.5000 1024.5850 1116.5000 1026.5850 ;
        RECT 1114.5000 1038.7750 1116.5000 1040.7750 ;
        RECT 1114.5000 1045.8700 1116.5000 1047.8700 ;
        RECT 1114.5000 1075.2500 1116.5000 1117.9000 ;
        RECT 1114.5000 1082.3450 1116.5000 1117.9000 ;
        RECT 1114.5000 1053.9650 1116.5000 1117.9000 ;
        RECT 1114.5000 1061.0600 1116.5000 1117.9000 ;
        RECT 1114.5000 1068.1550 1116.5000 1117.9000 ;
        RECT 1114.5000 1067.1550 1116.5000 1069.1550 ;
        RECT 1114.5000 1052.9650 1116.5000 1054.9650 ;
        RECT 1114.5000 1060.0600 1116.5000 1062.0600 ;
        RECT 1114.5000 1074.2500 1116.5000 1076.2500 ;
        RECT 1114.5000 1081.3450 1116.5000 1083.3450 ;
        RECT 1114.5000 1089.4400 1116.5000 1117.9000 ;
        RECT 1114.5000 1096.5350 1116.5000 1117.9000 ;
        RECT 1114.5000 1088.4400 1116.5000 1090.4400 ;
        RECT 1114.5000 1095.5350 1116.5000 1097.5350 ;
        RECT 1114.5000 1103.6300 1116.5000 1117.9000 ;
        RECT 1114.5000 1102.6300 1116.5000 1104.6300 ;
        RECT 1114.1000 138.2000 1116.1000 140.2000 ;
        RECT 1114.1000 47.0000 1116.1000 49.0000 ;
        RECT 1114.1000 60.2000 1116.1000 62.2000 ;
        RECT 1114.1000 53.0000 1116.1000 55.0000 ;
        RECT 1114.1000 67.2000 1116.1000 69.2000 ;
        RECT 1114.1000 74.4000 1116.1000 76.4000 ;
        RECT 1114.1000 81.4000 1116.1000 83.4000 ;
        RECT 1114.1000 95.6000 1116.1000 97.6000 ;
        RECT 1114.1000 88.6000 1116.1000 90.6000 ;
        RECT 1114.1000 102.8000 1116.1000 104.8000 ;
        RECT 1114.1000 109.8000 1116.1000 111.8000 ;
        RECT 1114.1000 117.0000 1116.1000 119.0000 ;
        RECT 1114.1000 131.2000 1116.1000 133.2000 ;
        RECT 1114.1000 124.0000 1116.1000 126.0000 ;
        RECT 1114.1000 209.2000 1116.1000 211.2000 ;
        RECT 1114.1000 173.6000 1116.1000 175.6000 ;
        RECT 1114.1000 145.4000 1116.1000 147.4000 ;
        RECT 1114.1000 152.4000 1116.1000 154.4000 ;
        RECT 1114.1000 159.4000 1116.1000 161.4000 ;
        RECT 1114.1000 166.6000 1116.1000 168.6000 ;
        RECT 1114.1000 180.8000 1116.1000 182.8000 ;
        RECT 1114.1000 187.8000 1116.1000 189.8000 ;
        RECT 1114.1000 195.0000 1116.1000 197.0000 ;
        RECT 1114.1000 202.0000 1116.1000 204.0000 ;
        RECT 1114.1000 244.6000 1116.1000 246.6000 ;
        RECT 1114.1000 216.2000 1116.1000 218.2000 ;
        RECT 1114.1000 223.4000 1116.1000 225.4000 ;
        RECT 1114.1000 230.4000 1116.1000 232.4000 ;
        RECT 1114.1000 237.6000 1116.1000 239.6000 ;
        RECT 1114.1000 251.8000 1116.1000 253.8000 ;
        RECT 1114.1000 258.8000 1116.1000 260.8000 ;
        RECT 1114.1000 266.4000 1116.1000 268.4000 ;
        RECT 1114.1000 273.6000 1116.1000 275.6000 ;
        RECT 1114.1000 287.2000 1116.1000 289.2000 ;
        RECT 1114.1000 280.8000 1116.1000 282.8000 ;
        RECT 1114.1000 294.4000 1116.1000 296.4000 ;
        RECT 1114.1000 301.4000 1116.1000 303.4000 ;
        RECT 1114.1000 308.4000 1116.1000 310.4000 ;
        RECT 1114.1000 322.6000 1116.1000 324.6000 ;
        RECT 1114.1000 315.6000 1116.1000 317.6000 ;
        RECT 1114.1000 329.8000 1116.1000 331.8000 ;
        RECT 1114.1000 336.8000 1116.1000 338.8000 ;
        RECT 1114.1000 344.0000 1116.1000 346.0000 ;
        RECT 1114.1000 358.2000 1116.1000 360.2000 ;
        RECT 1114.1000 351.0000 1116.1000 353.0000 ;
        RECT 1114.1000 365.2000 1116.1000 367.2000 ;
        RECT 1114.1000 373.6000 1116.1000 375.6000 ;
        RECT 1114.1000 400.8000 1116.1000 402.8000 ;
        RECT 1114.1000 386.6000 1116.1000 388.6000 ;
        RECT 1114.1000 393.8000 1116.1000 395.8000 ;
        RECT 1114.1000 407.8000 1116.1000 409.8000 ;
        RECT 1114.1000 415.0000 1116.1000 417.0000 ;
        RECT 1114.1000 436.2000 1116.1000 438.2000 ;
        RECT 1114.1000 422.0000 1116.1000 424.0000 ;
        RECT 1114.1000 429.2000 1116.1000 431.2000 ;
        RECT 1114.1000 443.2000 1116.1000 445.2000 ;
        RECT 1114.1000 450.4000 1116.1000 452.4000 ;
        RECT 1114.1000 471.6000 1116.1000 473.6000 ;
        RECT 1114.1000 457.4000 1116.1000 459.4000 ;
        RECT 1114.1000 464.6000 1116.1000 466.6000 ;
        RECT 1114.1000 478.8000 1116.1000 480.8000 ;
        RECT 1114.1000 485.8000 1116.1000 487.8000 ;
        RECT 1114.1000 507.2000 1116.1000 509.2000 ;
        RECT 1114.1000 493.0000 1116.1000 495.0000 ;
        RECT 1114.1000 500.0000 1116.1000 502.0000 ;
        RECT 1114.1000 514.8000 1116.1000 516.8000 ;
        RECT 1114.1000 522.0000 1116.1000 524.0000 ;
        RECT 1114.1000 528.4000 1116.1000 530.4000 ;
        RECT 1114.1000 535.6000 1116.1000 537.6000 ;
        RECT 1114.1000 549.8000 1116.1000 551.8000 ;
        RECT 1114.1000 542.6000 1116.1000 544.6000 ;
        RECT 1114.1000 556.8000 1116.1000 558.8000 ;
        RECT 1114.1000 698.8000 1116.1000 700.8000 ;
        RECT 1114.1000 564.0000 1116.1000 566.0000 ;
        RECT 1114.1000 571.0000 1116.1000 573.0000 ;
        RECT 1114.1000 585.2000 1116.1000 587.2000 ;
        RECT 1114.1000 578.2000 1116.1000 580.2000 ;
        RECT 1114.1000 592.2000 1116.1000 594.2000 ;
        RECT 1114.1000 599.4000 1116.1000 601.4000 ;
        RECT 1114.1000 606.4000 1116.1000 608.4000 ;
        RECT 1114.1000 620.6000 1116.1000 622.6000 ;
        RECT 1114.1000 613.6000 1116.1000 615.6000 ;
        RECT 1114.1000 627.8000 1116.1000 629.8000 ;
        RECT 1114.1000 663.2000 1116.1000 665.2000 ;
        RECT 1114.1000 634.8000 1116.1000 636.8000 ;
        RECT 1114.1000 642.0000 1116.1000 644.0000 ;
        RECT 1114.1000 656.2000 1116.1000 658.2000 ;
        RECT 1114.1000 649.0000 1116.1000 651.0000 ;
        RECT 1114.1000 670.4000 1116.1000 672.4000 ;
        RECT 1114.1000 677.4000 1116.1000 679.4000 ;
        RECT 1114.1000 684.6000 1116.1000 686.6000 ;
        RECT 1114.1000 691.6000 1116.1000 693.6000 ;
        RECT 1114.1000 705.8000 1116.1000 707.8000 ;
        RECT 1114.1000 713.0000 1116.1000 715.0000 ;
        RECT 1114.1000 720.0000 1116.1000 722.0000 ;
        RECT 1114.5000 721.0000 1116.5000 723.0000 ;
        RECT 2.0000 10.0000 4.0000 12.0000 ;
        RECT 106.5750 47.0000 108.5750 49.0000 ;
        RECT 106.5750 60.0700 108.5750 61.8350 ;
        RECT 1114.1000 279.6100 1118.0000 281.6100 ;
        RECT 1114.5000 17.0950 1118.0000 19.0950 ;
        RECT 1114.5000 10.0000 1118.0000 12.0000 ;
        RECT 1114.5000 24.1900 1118.0000 26.1900 ;
        RECT 1114.5000 31.2850 1118.0000 33.2850 ;
        RECT 1114.5000 38.3800 1118.0000 40.3800 ;
        RECT 1114.1000 45.4750 1118.0000 47.4750 ;
        RECT 1114.1000 59.6650 1118.0000 61.6650 ;
        RECT 1114.1000 52.5700 1118.0000 54.5700 ;
        RECT 1114.1000 66.7600 1118.0000 68.7600 ;
        RECT 1114.1000 73.8550 1118.0000 75.8550 ;
        RECT 1114.1000 80.9500 1118.0000 82.9500 ;
        RECT 1114.1000 95.1400 1118.0000 97.1400 ;
        RECT 1114.1000 88.0450 1118.0000 90.0450 ;
        RECT 1114.1000 102.2350 1118.0000 104.2350 ;
        RECT 1114.1000 109.3300 1118.0000 111.3300 ;
        RECT 1114.1000 116.4250 1118.0000 118.4250 ;
        RECT 1114.1000 130.6150 1118.0000 132.6150 ;
        RECT 1114.1000 123.5200 1118.0000 125.5200 ;
        RECT 1114.1000 137.7100 1118.0000 139.7100 ;
        RECT 1114.1000 208.6600 1118.0000 210.6600 ;
        RECT 1114.1000 173.1850 1118.0000 175.1850 ;
        RECT 1114.1000 144.8050 1118.0000 146.8050 ;
        RECT 1114.1000 151.9000 1118.0000 153.9000 ;
        RECT 1114.1000 166.0900 1118.0000 168.0900 ;
        RECT 1114.1000 158.9950 1118.0000 160.9950 ;
        RECT 1114.1000 180.2800 1118.0000 182.2800 ;
        RECT 1114.1000 187.3750 1118.0000 189.3750 ;
        RECT 1114.1000 194.4700 1118.0000 196.4700 ;
        RECT 1114.1000 201.5650 1118.0000 203.5650 ;
        RECT 1114.1000 244.1350 1118.0000 246.1350 ;
        RECT 1114.1000 215.7550 1118.0000 217.7550 ;
        RECT 1114.1000 222.8500 1118.0000 224.8500 ;
        RECT 1114.1000 229.9450 1118.0000 231.9450 ;
        RECT 1114.1000 237.0400 1118.0000 239.0400 ;
        RECT 1114.1000 251.2300 1118.0000 253.2300 ;
        RECT 1114.1000 258.3250 1118.0000 260.3250 ;
        RECT 1114.1000 265.4200 1118.0000 267.4200 ;
        RECT 1114.1000 272.5150 1118.0000 274.5150 ;
        RECT 1114.1000 286.7050 1118.0000 288.7050 ;
        RECT 1114.1000 293.8000 1118.0000 295.8000 ;
        RECT 1114.1000 300.8950 1118.0000 302.8950 ;
        RECT 1114.1000 307.9900 1118.0000 309.9900 ;
        RECT 1114.1000 322.1800 1118.0000 324.1800 ;
        RECT 1114.1000 315.0850 1118.0000 317.0850 ;
        RECT 1114.1000 329.2750 1118.0000 331.2750 ;
        RECT 1114.1000 336.3700 1118.0000 338.3700 ;
        RECT 1114.1000 343.4650 1118.0000 345.4650 ;
        RECT 1114.1000 357.6550 1118.0000 359.6550 ;
        RECT 1114.1000 350.5600 1118.0000 352.5600 ;
        RECT 1114.1000 364.7500 1118.0000 366.7500 ;
        RECT 1114.1000 371.8450 1118.0000 373.8450 ;
        RECT 1116.0000 378.9400 1118.0000 380.9400 ;
        RECT 1114.1000 393.1300 1118.0000 395.1300 ;
        RECT 1114.1000 386.0350 1118.0000 388.0350 ;
        RECT 1114.1000 400.2250 1118.0000 402.2250 ;
        RECT 1114.1000 407.3200 1118.0000 409.3200 ;
        RECT 1114.1000 414.4150 1118.0000 416.4150 ;
        RECT 1114.1000 435.7000 1118.0000 437.7000 ;
        RECT 1114.1000 428.6050 1118.0000 430.6050 ;
        RECT 1114.1000 421.5100 1118.0000 423.5100 ;
        RECT 1114.1000 442.7950 1118.0000 444.7950 ;
        RECT 1114.1000 449.8900 1118.0000 451.8900 ;
        RECT 1114.1000 471.1750 1118.0000 473.1750 ;
        RECT 1114.1000 456.9850 1118.0000 458.9850 ;
        RECT 1114.1000 464.0800 1118.0000 466.0800 ;
        RECT 1114.1000 478.2700 1118.0000 480.2700 ;
        RECT 1114.1000 485.3650 1118.0000 487.3650 ;
        RECT 1114.1000 506.6500 1118.0000 508.6500 ;
        RECT 1114.1000 492.4600 1118.0000 494.4600 ;
        RECT 1114.1000 499.5550 1118.0000 501.5550 ;
        RECT 1114.1000 513.7450 1118.0000 515.7450 ;
        RECT 1114.1000 520.8400 1118.0000 522.8400 ;
        RECT 1114.1000 542.1250 1118.0000 544.1250 ;
        RECT 1114.1000 527.9350 1118.0000 529.9350 ;
        RECT 1114.1000 535.0300 1118.0000 537.0300 ;
        RECT 1114.1000 549.2200 1118.0000 551.2200 ;
        RECT 1114.1000 556.3150 1118.0000 558.3150 ;
        RECT 2.0000 804.6400 4.0000 806.6400 ;
        RECT 2.0000 790.4500 4.0000 792.4500 ;
        RECT 2.0000 797.5450 4.0000 799.5450 ;
        RECT 2.0000 811.7350 4.0000 813.7350 ;
        RECT 2.0000 818.8300 4.0000 820.8300 ;
        RECT 2.0000 825.9250 4.0000 827.9250 ;
        RECT 2.0000 833.0200 4.0000 835.0200 ;
        RECT 327.9650 678.1650 329.9650 679.3350 ;
        RECT 327.9650 691.5250 329.9650 693.0000 ;
        RECT 410.1500 708.1650 412.1500 709.8100 ;
        RECT 410.1500 721.0000 412.1500 723.0000 ;
        RECT 2.0000 847.2100 4.0000 849.2100 ;
        RECT 2.0000 840.1150 4.0000 842.1150 ;
        RECT 2.0000 854.3050 4.0000 856.3050 ;
        RECT 2.0000 861.4000 4.0000 863.4000 ;
        RECT 2.0000 868.4950 4.0000 870.4950 ;
        RECT 2.0000 882.6850 4.0000 884.6850 ;
        RECT 2.0000 875.5900 4.0000 877.5900 ;
        RECT 2.0000 889.7800 4.0000 891.7800 ;
        RECT 2.0000 896.8750 4.0000 898.8750 ;
        RECT 2.0000 903.9700 4.0000 905.9700 ;
        RECT 2.0000 918.1600 4.0000 920.1600 ;
        RECT 2.0000 911.0650 4.0000 913.0650 ;
        RECT 2.0000 925.2550 4.0000 927.2550 ;
        RECT 2.0000 932.3500 4.0000 934.3500 ;
        RECT 2.0000 939.4450 4.0000 941.4450 ;
        RECT 2.0000 960.7300 4.0000 962.7300 ;
        RECT 2.0000 953.6350 4.0000 955.6350 ;
        RECT 2.0000 946.5400 4.0000 948.5400 ;
        RECT 2.0000 967.8250 4.0000 969.8250 ;
        RECT 2.0000 974.9200 4.0000 976.9200 ;
        RECT 2.0000 996.2050 4.0000 998.2050 ;
        RECT 2.0000 982.0150 4.0000 984.0150 ;
        RECT 2.0000 989.1100 4.0000 991.1100 ;
        RECT 2.0000 1003.3000 4.0000 1005.3000 ;
        RECT 1114.1000 698.2150 1118.0000 700.2150 ;
        RECT 1114.1000 563.4100 1118.0000 565.4100 ;
        RECT 1114.1000 570.5050 1118.0000 572.5050 ;
        RECT 1114.1000 584.6950 1118.0000 586.6950 ;
        RECT 1114.1000 577.6000 1118.0000 579.6000 ;
        RECT 1114.1000 591.7900 1118.0000 593.7900 ;
        RECT 1114.1000 598.8850 1118.0000 600.8850 ;
        RECT 1114.1000 605.9800 1118.0000 607.9800 ;
        RECT 1114.1000 620.1700 1118.0000 622.1700 ;
        RECT 1114.1000 613.0750 1118.0000 615.0750 ;
        RECT 1114.1000 627.2650 1118.0000 629.2650 ;
        RECT 1114.1000 634.3600 1118.0000 636.3600 ;
        RECT 1114.1000 641.4550 1118.0000 643.4550 ;
        RECT 1114.1000 655.6450 1118.0000 657.6450 ;
        RECT 1114.1000 648.5500 1118.0000 650.5500 ;
        RECT 1114.1000 662.7400 1118.0000 664.7400 ;
        RECT 1114.1000 669.8350 1118.0000 671.8350 ;
        RECT 1114.1000 676.9300 1118.0000 678.9300 ;
        RECT 1114.1000 691.1200 1118.0000 693.1200 ;
        RECT 1114.1000 684.0250 1118.0000 686.0250 ;
        RECT 1114.5000 769.1650 1118.0000 771.1650 ;
        RECT 1114.5000 733.6900 1118.0000 735.6900 ;
        RECT 1114.1000 705.3100 1118.0000 707.3100 ;
        RECT 1114.1000 712.4050 1118.0000 714.4050 ;
        RECT 1114.1000 719.5000 1118.0000 721.5000 ;
        RECT 1114.5000 726.5950 1118.0000 728.5950 ;
        RECT 1114.5000 740.7850 1118.0000 742.7850 ;
        RECT 1114.5000 747.8800 1118.0000 749.8800 ;
        RECT 1114.5000 754.9750 1118.0000 756.9750 ;
        RECT 1114.5000 762.0700 1118.0000 764.0700 ;
        RECT 1116.0000 804.6400 1118.0000 806.6400 ;
        RECT 1114.5000 776.2600 1118.0000 778.2600 ;
        RECT 1114.5000 783.3550 1118.0000 785.3550 ;
        RECT 1116.0000 790.4500 1118.0000 792.4500 ;
        RECT 1114.7150 791.0350 1115.1250 791.3650 ;
        RECT 1116.0000 797.5450 1118.0000 799.5450 ;
        RECT 1114.7150 798.2350 1115.1250 798.5650 ;
        RECT 1114.7150 805.4350 1115.1250 805.7650 ;
        RECT 1114.7150 812.6350 1115.1250 812.9650 ;
        RECT 1116.0000 811.7350 1118.0000 813.7350 ;
        RECT 1116.0000 818.8300 1118.0000 820.8300 ;
        RECT 1114.7150 819.8350 1115.1250 820.1650 ;
        RECT 1114.7150 827.0350 1115.1250 827.3650 ;
        RECT 1116.0000 825.9250 1118.0000 827.9250 ;
        RECT 1116.0000 833.0200 1118.0000 835.0200 ;
        RECT 1114.7150 834.2350 1115.1250 834.5650 ;
        RECT 1116.0000 847.2100 1118.0000 849.2100 ;
        RECT 1114.7150 848.6350 1115.1250 848.9650 ;
        RECT 1116.0000 840.1150 1118.0000 842.1150 ;
        RECT 1114.7150 841.4350 1115.1250 841.7650 ;
        RECT 1116.0000 854.3050 1118.0000 856.3050 ;
        RECT 1114.7150 855.8350 1115.1250 856.1650 ;
        RECT 1116.0000 861.4000 1118.0000 863.4000 ;
        RECT 1114.7150 863.0350 1115.1250 863.3650 ;
        RECT 1116.0000 868.4950 1118.0000 870.4950 ;
        RECT 1116.0000 882.6850 1118.0000 884.6850 ;
        RECT 1116.0000 875.5900 1118.0000 877.5900 ;
        RECT 1116.0000 889.7800 1118.0000 891.7800 ;
        RECT 1116.0000 896.8750 1118.0000 898.8750 ;
        RECT 1116.0000 903.9700 1118.0000 905.9700 ;
        RECT 1116.0000 918.1600 1118.0000 920.1600 ;
        RECT 1116.0000 911.0650 1118.0000 913.0650 ;
        RECT 1116.0000 925.2550 1118.0000 927.2550 ;
        RECT 1116.0000 932.3500 1118.0000 934.3500 ;
        RECT 1116.0000 939.4450 1118.0000 941.4450 ;
        RECT 1116.0000 960.7300 1118.0000 962.7300 ;
        RECT 1116.0000 953.6350 1118.0000 955.6350 ;
        RECT 1116.0000 946.5400 1118.0000 948.5400 ;
        RECT 1116.0000 967.8250 1118.0000 969.8250 ;
        RECT 1116.0000 974.9200 1118.0000 976.9200 ;
        RECT 1116.0000 996.2050 1118.0000 998.2050 ;
        RECT 1116.0000 982.0150 1118.0000 984.0150 ;
        RECT 1114.7150 996.2350 1115.1250 996.5650 ;
        RECT 1116.0000 989.1100 1118.0000 991.1100 ;
        RECT 1116.0000 1003.3000 1118.0000 1005.3000 ;
        RECT 1114.7150 1003.4350 1115.1250 1003.7650 ;
        RECT 1114.5000 1010.3950 1118.0000 1012.3950 ;
        RECT 1114.5000 1031.6800 1118.0000 1033.6800 ;
        RECT 1114.5000 1017.4900 1118.0000 1019.4900 ;
        RECT 1114.5000 1024.5850 1118.0000 1026.5850 ;
        RECT 1114.5000 1038.7750 1118.0000 1040.7750 ;
        RECT 1114.5000 1045.8700 1118.0000 1047.8700 ;
        RECT 1114.5000 1067.1550 1118.0000 1069.1550 ;
        RECT 1114.5000 1052.9650 1118.0000 1054.9650 ;
        RECT 1114.5000 1060.0600 1118.0000 1062.0600 ;
        RECT 1114.5000 1074.2500 1118.0000 1076.2500 ;
        RECT 1114.5000 1081.3450 1118.0000 1083.3450 ;
        RECT 1114.5000 1088.4400 1118.0000 1090.4400 ;
        RECT 1114.5000 1095.5350 1118.0000 1097.5350 ;
        RECT 1114.5000 1102.6300 1118.0000 1104.6300 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'sram_w16_64b'
    PORT
      LAYER M4 ;
        RECT 327.9650 329.8350 329.9650 330.1650 ;
        RECT 319.4500 329.8350 321.4500 330.1650 ;
        RECT 310.9350 329.8350 312.9350 330.1650 ;
        RECT 293.9050 329.8350 295.9050 330.1650 ;
        RECT 276.8750 329.8350 278.8750 330.1650 ;
        RECT 268.3600 329.8350 270.3600 330.1650 ;
        RECT 285.3900 329.8350 287.3900 330.1650 ;
        RECT 302.4200 329.8350 304.4200 330.1650 ;
        RECT 259.8450 329.8350 261.8450 330.1650 ;
        RECT 251.3300 329.8350 253.3300 330.1650 ;
        RECT 242.8150 329.8350 244.8150 330.1650 ;
        RECT 234.3000 329.8350 236.3000 330.1650 ;
        RECT 225.7850 329.8350 227.7850 330.1650 ;
        RECT 217.2700 329.8350 219.2700 330.1650 ;
        RECT 208.7550 329.8350 210.7550 330.1650 ;
        RECT 200.2400 329.8350 202.2400 330.1650 ;
        RECT 191.7250 329.8350 193.7250 330.1650 ;
        RECT 183.2100 329.8350 185.2100 330.1650 ;
        RECT 174.6950 329.8350 176.6950 330.1650 ;
        RECT 166.1800 329.8350 168.1800 330.1650 ;
        RECT 140.6350 329.8350 142.6350 330.1650 ;
        RECT 149.1500 329.8350 151.1500 330.1650 ;
        RECT 132.1200 329.8350 134.1200 330.1650 ;
        RECT 123.6050 329.8350 125.6050 330.1650 ;
        RECT 157.6650 329.8350 159.6650 330.1650 ;
        RECT 115.0900 329.8350 117.0900 330.1650 ;
        RECT 106.5750 329.8350 108.5750 330.1650 ;
        RECT 98.0600 329.8350 100.0600 330.1650 ;
        RECT 89.5450 329.8350 91.5450 330.1650 ;
        RECT 81.0300 329.8350 83.0300 330.1650 ;
        RECT 72.5150 329.8350 74.5150 330.1650 ;
        RECT 64.0000 329.8350 66.0000 330.1650 ;
        RECT 327.9650 59.8350 329.9650 60.1650 ;
        RECT 319.4500 59.8350 321.4500 60.1650 ;
        RECT 310.9350 59.8350 312.9350 60.1650 ;
        RECT 293.9050 59.8350 295.9050 60.1650 ;
        RECT 276.8750 59.8350 278.8750 60.1650 ;
        RECT 268.3600 59.8350 270.3600 60.1650 ;
        RECT 285.3900 59.8350 287.3900 60.1650 ;
        RECT 302.4200 59.8350 304.4200 60.1650 ;
        RECT 259.8450 59.8350 261.8450 60.1650 ;
        RECT 251.3300 59.8350 253.3300 60.1650 ;
        RECT 242.8150 59.8350 244.8150 60.1650 ;
        RECT 234.3000 59.8350 236.3000 60.1650 ;
        RECT 225.7850 59.8350 227.7850 60.1650 ;
        RECT 217.2700 59.8350 219.2700 60.1650 ;
        RECT 208.7550 59.8350 210.7550 60.1650 ;
        RECT 200.2400 59.8350 202.2400 60.1650 ;
        RECT 191.7250 59.8350 193.7250 60.1650 ;
        RECT 183.2100 59.8350 185.2100 60.1650 ;
        RECT 174.6950 59.8350 176.6950 60.1650 ;
        RECT 166.1800 59.8350 168.1800 60.1650 ;
        RECT 140.6350 59.8350 142.6350 60.1650 ;
        RECT 149.1500 59.8350 151.1500 60.1650 ;
        RECT 132.1200 59.8350 134.1200 60.1650 ;
        RECT 123.6050 59.8350 125.6050 60.1650 ;
        RECT 157.6650 59.8350 159.6650 60.1650 ;
        RECT 115.0900 59.8350 117.0900 60.1650 ;
        RECT 106.5750 59.8350 108.5750 60.1650 ;
        RECT 98.0600 59.8350 100.0600 60.1650 ;
        RECT 89.5450 59.8350 91.5450 60.1650 ;
        RECT 81.0300 59.8350 83.0300 60.1650 ;
        RECT 72.5150 59.8350 74.5150 60.1650 ;
        RECT 64.0000 59.8350 66.0000 60.1650 ;
        RECT 310.9350 60.0000 312.9350 330.0000 ;
        RECT 319.4500 60.0000 321.4500 330.0000 ;
        RECT 327.9650 60.0000 329.9650 330.0000 ;
        RECT 293.9050 60.0000 295.9050 330.0000 ;
        RECT 268.3600 60.0000 270.3600 330.0000 ;
        RECT 276.8750 60.0000 278.8750 330.0000 ;
        RECT 285.3900 60.0000 287.3900 330.0000 ;
        RECT 302.4200 60.0000 304.4200 330.0000 ;
        RECT 251.3300 60.0000 253.3300 330.0000 ;
        RECT 259.8450 60.0000 261.8450 330.0000 ;
        RECT 234.3000 60.0000 236.3000 330.0000 ;
        RECT 242.8150 60.0000 244.8150 330.0000 ;
        RECT 217.2700 60.0000 219.2700 330.0000 ;
        RECT 225.7850 60.0000 227.7850 330.0000 ;
        RECT 200.2400 60.0000 202.2400 330.0000 ;
        RECT 208.7550 60.0000 210.7550 330.0000 ;
        RECT 191.7250 60.0000 193.7250 330.0000 ;
        RECT 183.2100 60.0000 185.2100 330.0000 ;
        RECT 166.1800 60.0000 168.1800 330.0000 ;
        RECT 174.6950 60.0000 176.6950 330.0000 ;
        RECT 140.6350 60.0000 142.6350 330.0000 ;
        RECT 149.1500 60.0000 151.1500 330.0000 ;
        RECT 123.6050 60.0000 125.6050 330.0000 ;
        RECT 132.1200 60.0000 134.1200 330.0000 ;
        RECT 157.6650 60.0000 159.6650 330.0000 ;
        RECT 106.5750 60.0000 108.5750 330.0000 ;
        RECT 115.0900 60.0000 117.0900 330.0000 ;
        RECT 89.5450 60.0000 91.5450 330.0000 ;
        RECT 98.0600 60.0000 100.0600 330.0000 ;
        RECT 81.0300 60.0000 83.0300 330.0000 ;
        RECT 72.5150 60.0000 74.5150 330.0000 ;
        RECT 64.0000 60.0000 66.0000 330.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16_64b'


# P/G pin shape extracted from block 'sram_w16_64b'
    PORT
      LAYER M4 ;
        RECT 327.9650 679.8350 329.9650 680.1650 ;
        RECT 319.4500 679.8350 321.4500 680.1650 ;
        RECT 310.9350 679.8350 312.9350 680.1650 ;
        RECT 293.9050 679.8350 295.9050 680.1650 ;
        RECT 276.8750 679.8350 278.8750 680.1650 ;
        RECT 268.3600 679.8350 270.3600 680.1650 ;
        RECT 285.3900 679.8350 287.3900 680.1650 ;
        RECT 302.4200 679.8350 304.4200 680.1650 ;
        RECT 259.8450 679.8350 261.8450 680.1650 ;
        RECT 251.3300 679.8350 253.3300 680.1650 ;
        RECT 242.8150 679.8350 244.8150 680.1650 ;
        RECT 234.3000 679.8350 236.3000 680.1650 ;
        RECT 225.7850 679.8350 227.7850 680.1650 ;
        RECT 217.2700 679.8350 219.2700 680.1650 ;
        RECT 208.7550 679.8350 210.7550 680.1650 ;
        RECT 200.2400 679.8350 202.2400 680.1650 ;
        RECT 191.7250 679.8350 193.7250 680.1650 ;
        RECT 183.2100 679.8350 185.2100 680.1650 ;
        RECT 174.6950 679.8350 176.6950 680.1650 ;
        RECT 166.1800 679.8350 168.1800 680.1650 ;
        RECT 140.6350 679.8350 142.6350 680.1650 ;
        RECT 149.1500 679.8350 151.1500 680.1650 ;
        RECT 132.1200 679.8350 134.1200 680.1650 ;
        RECT 123.6050 679.8350 125.6050 680.1650 ;
        RECT 157.6650 679.8350 159.6650 680.1650 ;
        RECT 115.0900 679.8350 117.0900 680.1650 ;
        RECT 106.5750 679.8350 108.5750 680.1650 ;
        RECT 98.0600 679.8350 100.0600 680.1650 ;
        RECT 89.5450 679.8350 91.5450 680.1650 ;
        RECT 81.0300 679.8350 83.0300 680.1650 ;
        RECT 72.5150 679.8350 74.5150 680.1650 ;
        RECT 64.0000 679.8350 66.0000 680.1650 ;
        RECT 327.9650 409.8350 329.9650 410.1650 ;
        RECT 319.4500 409.8350 321.4500 410.1650 ;
        RECT 310.9350 409.8350 312.9350 410.1650 ;
        RECT 293.9050 409.8350 295.9050 410.1650 ;
        RECT 276.8750 409.8350 278.8750 410.1650 ;
        RECT 268.3600 409.8350 270.3600 410.1650 ;
        RECT 285.3900 409.8350 287.3900 410.1650 ;
        RECT 302.4200 409.8350 304.4200 410.1650 ;
        RECT 259.8450 409.8350 261.8450 410.1650 ;
        RECT 251.3300 409.8350 253.3300 410.1650 ;
        RECT 242.8150 409.8350 244.8150 410.1650 ;
        RECT 234.3000 409.8350 236.3000 410.1650 ;
        RECT 225.7850 409.8350 227.7850 410.1650 ;
        RECT 217.2700 409.8350 219.2700 410.1650 ;
        RECT 208.7550 409.8350 210.7550 410.1650 ;
        RECT 200.2400 409.8350 202.2400 410.1650 ;
        RECT 191.7250 409.8350 193.7250 410.1650 ;
        RECT 183.2100 409.8350 185.2100 410.1650 ;
        RECT 174.6950 409.8350 176.6950 410.1650 ;
        RECT 166.1800 409.8350 168.1800 410.1650 ;
        RECT 140.6350 409.8350 142.6350 410.1650 ;
        RECT 149.1500 409.8350 151.1500 410.1650 ;
        RECT 132.1200 409.8350 134.1200 410.1650 ;
        RECT 123.6050 409.8350 125.6050 410.1650 ;
        RECT 157.6650 409.8350 159.6650 410.1650 ;
        RECT 115.0900 409.8350 117.0900 410.1650 ;
        RECT 106.5750 409.8350 108.5750 410.1650 ;
        RECT 98.0600 409.8350 100.0600 410.1650 ;
        RECT 89.5450 409.8350 91.5450 410.1650 ;
        RECT 81.0300 409.8350 83.0300 410.1650 ;
        RECT 72.5150 409.8350 74.5150 410.1650 ;
        RECT 64.0000 409.8350 66.0000 410.1650 ;
        RECT 310.9350 410.0000 312.9350 680.0000 ;
        RECT 319.4500 410.0000 321.4500 680.0000 ;
        RECT 327.9650 410.0000 329.9650 680.0000 ;
        RECT 293.9050 410.0000 295.9050 680.0000 ;
        RECT 268.3600 410.0000 270.3600 680.0000 ;
        RECT 276.8750 410.0000 278.8750 680.0000 ;
        RECT 285.3900 410.0000 287.3900 680.0000 ;
        RECT 302.4200 410.0000 304.4200 680.0000 ;
        RECT 251.3300 410.0000 253.3300 680.0000 ;
        RECT 259.8450 410.0000 261.8450 680.0000 ;
        RECT 234.3000 410.0000 236.3000 680.0000 ;
        RECT 242.8150 410.0000 244.8150 680.0000 ;
        RECT 217.2700 410.0000 219.2700 680.0000 ;
        RECT 225.7850 410.0000 227.7850 680.0000 ;
        RECT 200.2400 410.0000 202.2400 680.0000 ;
        RECT 208.7550 410.0000 210.7550 680.0000 ;
        RECT 191.7250 410.0000 193.7250 680.0000 ;
        RECT 183.2100 410.0000 185.2100 680.0000 ;
        RECT 166.1800 410.0000 168.1800 680.0000 ;
        RECT 174.6950 410.0000 176.6950 680.0000 ;
        RECT 140.6350 410.0000 142.6350 680.0000 ;
        RECT 149.1500 410.0000 151.1500 680.0000 ;
        RECT 123.6050 410.0000 125.6050 680.0000 ;
        RECT 132.1200 410.0000 134.1200 680.0000 ;
        RECT 157.6650 410.0000 159.6650 680.0000 ;
        RECT 106.5750 410.0000 108.5750 680.0000 ;
        RECT 115.0900 410.0000 117.0900 680.0000 ;
        RECT 89.5450 410.0000 91.5450 680.0000 ;
        RECT 98.0600 410.0000 100.0600 680.0000 ;
        RECT 81.0300 410.0000 83.0300 680.0000 ;
        RECT 72.5150 410.0000 74.5150 680.0000 ;
        RECT 64.0000 410.0000 66.0000 680.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16_64b'


# P/G pin shape extracted from block 'sram_w16_160b'
    PORT
      LAYER M4 ;
        RECT 418.3000 709.8350 420.3000 710.1650 ;
        RECT 410.1500 709.8350 412.1500 710.1650 ;
        RECT 434.6000 709.8350 436.6000 710.1650 ;
        RECT 426.4500 709.8350 428.4500 710.1650 ;
        RECT 459.0500 709.8350 461.0500 710.1650 ;
        RECT 450.9000 709.8350 452.9000 710.1650 ;
        RECT 442.7500 709.8350 444.7500 710.1650 ;
        RECT 475.3500 709.8350 477.3500 710.1650 ;
        RECT 467.2000 709.8350 469.2000 710.1650 ;
        RECT 499.8000 709.8350 501.8000 710.1650 ;
        RECT 491.6500 709.8350 493.6500 710.1650 ;
        RECT 516.1000 709.8350 518.1000 710.1650 ;
        RECT 507.9500 709.8350 509.9500 710.1650 ;
        RECT 540.5500 709.8350 542.5500 710.1650 ;
        RECT 532.4000 709.8350 534.4000 710.1650 ;
        RECT 565.0000 709.8350 567.0000 710.1650 ;
        RECT 556.8500 709.8350 558.8500 710.1650 ;
        RECT 548.7000 709.8350 550.7000 710.1650 ;
        RECT 524.2500 709.8350 526.2500 710.1650 ;
        RECT 483.5000 709.8350 485.5000 710.1650 ;
        RECT 581.3000 709.8350 583.3000 710.1650 ;
        RECT 573.1500 709.8350 575.1500 710.1650 ;
        RECT 605.7500 709.8350 607.7500 710.1650 ;
        RECT 597.6000 709.8350 599.6000 710.1650 ;
        RECT 589.4500 709.8350 591.4500 710.1650 ;
        RECT 622.0500 709.8350 624.0500 710.1650 ;
        RECT 613.9000 709.8350 615.9000 710.1650 ;
        RECT 646.5000 709.8350 648.5000 710.1650 ;
        RECT 638.3500 709.8350 640.3500 710.1650 ;
        RECT 630.2000 709.8350 632.2000 710.1650 ;
        RECT 662.8000 709.8350 664.8000 710.1650 ;
        RECT 654.6500 709.8350 656.6500 710.1650 ;
        RECT 687.2500 709.8350 689.2500 710.1650 ;
        RECT 679.1000 709.8350 681.1000 710.1650 ;
        RECT 670.9500 709.8350 672.9500 710.1650 ;
        RECT 711.7000 709.8350 713.7000 710.1650 ;
        RECT 703.5500 709.8350 705.5500 710.1650 ;
        RECT 695.4000 709.8350 697.4000 710.1650 ;
        RECT 728.0000 709.8350 730.0000 710.1650 ;
        RECT 719.8500 709.8350 721.8500 710.1650 ;
        RECT 752.4500 709.8350 754.4500 710.1650 ;
        RECT 744.3000 709.8350 746.3000 710.1650 ;
        RECT 736.1500 709.8350 738.1500 710.1650 ;
        RECT 768.7500 709.8350 770.7500 710.1650 ;
        RECT 760.6000 709.8350 762.6000 710.1650 ;
        RECT 793.2000 709.8350 795.2000 710.1650 ;
        RECT 785.0500 709.8350 787.0500 710.1650 ;
        RECT 776.9000 709.8350 778.9000 710.1650 ;
        RECT 809.5000 709.8350 811.5000 710.1650 ;
        RECT 801.3500 709.8350 803.3500 710.1650 ;
        RECT 833.9500 709.8350 835.9500 710.1650 ;
        RECT 825.8000 709.8350 827.8000 710.1650 ;
        RECT 858.4000 709.8350 860.4000 710.1650 ;
        RECT 850.2500 709.8350 852.2500 710.1650 ;
        RECT 842.1000 709.8350 844.1000 710.1650 ;
        RECT 874.7000 709.8350 876.7000 710.1650 ;
        RECT 866.5500 709.8350 868.5500 710.1650 ;
        RECT 899.1500 709.8350 901.1500 710.1650 ;
        RECT 891.0000 709.8350 893.0000 710.1650 ;
        RECT 882.8500 709.8350 884.8500 710.1650 ;
        RECT 817.6500 709.8350 819.6500 710.1650 ;
        RECT 915.4500 709.8350 917.4500 710.1650 ;
        RECT 907.3000 709.8350 909.3000 710.1650 ;
        RECT 939.9000 709.8350 941.9000 710.1650 ;
        RECT 931.7500 709.8350 933.7500 710.1650 ;
        RECT 923.6000 709.8350 925.6000 710.1650 ;
        RECT 956.2000 709.8350 958.2000 710.1650 ;
        RECT 948.0500 709.8350 950.0500 710.1650 ;
        RECT 980.6500 709.8350 982.6500 710.1650 ;
        RECT 972.5000 709.8350 974.5000 710.1650 ;
        RECT 964.3500 709.8350 966.3500 710.1650 ;
        RECT 1005.1000 709.8350 1007.1000 710.1650 ;
        RECT 996.9500 709.8350 998.9500 710.1650 ;
        RECT 988.8000 709.8350 990.8000 710.1650 ;
        RECT 1021.4000 709.8350 1023.4000 710.1650 ;
        RECT 1013.2500 709.8350 1015.2500 710.1650 ;
        RECT 1045.8500 709.8350 1047.8500 710.1650 ;
        RECT 1037.7000 709.8350 1039.7000 710.1650 ;
        RECT 1029.5500 709.8350 1031.5500 710.1650 ;
        RECT 1054.0000 709.8350 1056.0000 710.1650 ;
        RECT 410.1500 60.0000 412.1500 710.0000 ;
        RECT 418.3000 60.0000 420.3000 710.0000 ;
        RECT 426.4500 60.0000 428.4500 710.0000 ;
        RECT 434.6000 60.0000 436.6000 710.0000 ;
        RECT 442.7500 60.0000 444.7500 710.0000 ;
        RECT 450.9000 60.0000 452.9000 710.0000 ;
        RECT 459.0500 60.0000 461.0500 710.0000 ;
        RECT 467.2000 60.0000 469.2000 710.0000 ;
        RECT 475.3500 60.0000 477.3500 710.0000 ;
        RECT 565.0000 60.0000 567.0000 710.0000 ;
        RECT 556.8500 60.0000 558.8500 710.0000 ;
        RECT 548.7000 60.0000 550.7000 710.0000 ;
        RECT 540.5500 60.0000 542.5500 710.0000 ;
        RECT 532.4000 60.0000 534.4000 710.0000 ;
        RECT 524.2500 60.0000 526.2500 710.0000 ;
        RECT 516.1000 60.0000 518.1000 710.0000 ;
        RECT 507.9500 60.0000 509.9500 710.0000 ;
        RECT 499.8000 60.0000 501.8000 710.0000 ;
        RECT 491.6500 60.0000 493.6500 710.0000 ;
        RECT 483.5000 60.0000 485.5000 710.0000 ;
        RECT 573.1500 60.0000 575.1500 710.0000 ;
        RECT 581.3000 60.0000 583.3000 710.0000 ;
        RECT 589.4500 60.0000 591.4500 710.0000 ;
        RECT 597.6000 60.0000 599.6000 710.0000 ;
        RECT 605.7500 60.0000 607.7500 710.0000 ;
        RECT 613.9000 60.0000 615.9000 710.0000 ;
        RECT 622.0500 60.0000 624.0500 710.0000 ;
        RECT 630.2000 60.0000 632.2000 710.0000 ;
        RECT 638.3500 60.0000 640.3500 710.0000 ;
        RECT 646.5000 60.0000 648.5000 710.0000 ;
        RECT 654.6500 60.0000 656.6500 710.0000 ;
        RECT 728.0000 60.0000 730.0000 710.0000 ;
        RECT 719.8500 60.0000 721.8500 710.0000 ;
        RECT 711.7000 60.0000 713.7000 710.0000 ;
        RECT 703.5500 60.0000 705.5500 710.0000 ;
        RECT 695.4000 60.0000 697.4000 710.0000 ;
        RECT 687.2500 60.0000 689.2500 710.0000 ;
        RECT 679.1000 60.0000 681.1000 710.0000 ;
        RECT 670.9500 60.0000 672.9500 710.0000 ;
        RECT 662.8000 60.0000 664.8000 710.0000 ;
        RECT 736.1500 60.0000 738.1500 710.0000 ;
        RECT 744.3000 60.0000 746.3000 710.0000 ;
        RECT 752.4500 60.0000 754.4500 710.0000 ;
        RECT 760.6000 60.0000 762.6000 710.0000 ;
        RECT 768.7500 60.0000 770.7500 710.0000 ;
        RECT 776.9000 60.0000 778.9000 710.0000 ;
        RECT 785.0500 60.0000 787.0500 710.0000 ;
        RECT 793.2000 60.0000 795.2000 710.0000 ;
        RECT 801.3500 60.0000 803.3500 710.0000 ;
        RECT 809.5000 60.0000 811.5000 710.0000 ;
        RECT 899.1500 60.0000 901.1500 710.0000 ;
        RECT 891.0000 60.0000 893.0000 710.0000 ;
        RECT 882.8500 60.0000 884.8500 710.0000 ;
        RECT 874.7000 60.0000 876.7000 710.0000 ;
        RECT 866.5500 60.0000 868.5500 710.0000 ;
        RECT 858.4000 60.0000 860.4000 710.0000 ;
        RECT 850.2500 60.0000 852.2500 710.0000 ;
        RECT 842.1000 60.0000 844.1000 710.0000 ;
        RECT 833.9500 60.0000 835.9500 710.0000 ;
        RECT 825.8000 60.0000 827.8000 710.0000 ;
        RECT 817.6500 60.0000 819.6500 710.0000 ;
        RECT 907.3000 60.0000 909.3000 710.0000 ;
        RECT 915.4500 60.0000 917.4500 710.0000 ;
        RECT 923.6000 60.0000 925.6000 710.0000 ;
        RECT 931.7500 60.0000 933.7500 710.0000 ;
        RECT 939.9000 60.0000 941.9000 710.0000 ;
        RECT 948.0500 60.0000 950.0500 710.0000 ;
        RECT 956.2000 60.0000 958.2000 710.0000 ;
        RECT 964.3500 60.0000 966.3500 710.0000 ;
        RECT 972.5000 60.0000 974.5000 710.0000 ;
        RECT 980.6500 60.0000 982.6500 710.0000 ;
        RECT 1054.0000 60.0000 1056.0000 710.0000 ;
        RECT 1045.8500 60.0000 1047.8500 710.0000 ;
        RECT 1037.7000 60.0000 1039.7000 710.0000 ;
        RECT 1029.5500 60.0000 1031.5500 710.0000 ;
        RECT 1021.4000 60.0000 1023.4000 710.0000 ;
        RECT 1013.2500 60.0000 1015.2500 710.0000 ;
        RECT 1005.1000 60.0000 1007.1000 710.0000 ;
        RECT 996.9500 60.0000 998.9500 710.0000 ;
        RECT 988.8000 60.0000 990.8000 710.0000 ;
    END
# end of P/G pin shape extracted from block 'sram_w16_160b'

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1120.0000 1120.0000 ;
    LAYER M2 ;
      RECT 724.0500 1119.3800 1120.0000 1120.0000 ;
      RECT 720.0500 1119.3800 723.7500 1120.0000 ;
      RECT 716.0500 1119.3800 719.7500 1120.0000 ;
      RECT 712.0500 1119.3800 715.7500 1120.0000 ;
      RECT 708.0500 1119.3800 711.7500 1120.0000 ;
      RECT 704.0500 1119.3800 707.7500 1120.0000 ;
      RECT 700.0500 1119.3800 703.7500 1120.0000 ;
      RECT 696.0500 1119.3800 699.7500 1120.0000 ;
      RECT 692.0500 1119.3800 695.7500 1120.0000 ;
      RECT 688.0500 1119.3800 691.7500 1120.0000 ;
      RECT 684.0500 1119.3800 687.7500 1120.0000 ;
      RECT 680.0500 1119.3800 683.7500 1120.0000 ;
      RECT 676.0500 1119.3800 679.7500 1120.0000 ;
      RECT 672.0500 1119.3800 675.7500 1120.0000 ;
      RECT 668.0500 1119.3800 671.7500 1120.0000 ;
      RECT 664.0500 1119.3800 667.7500 1120.0000 ;
      RECT 660.0500 1119.3800 663.7500 1120.0000 ;
      RECT 656.0500 1119.3800 659.7500 1120.0000 ;
      RECT 652.0500 1119.3800 655.7500 1120.0000 ;
      RECT 648.0500 1119.3800 651.7500 1120.0000 ;
      RECT 644.0500 1119.3800 647.7500 1120.0000 ;
      RECT 640.0500 1119.3800 643.7500 1120.0000 ;
      RECT 636.0500 1119.3800 639.7500 1120.0000 ;
      RECT 632.0500 1119.3800 635.7500 1120.0000 ;
      RECT 628.0500 1119.3800 631.7500 1120.0000 ;
      RECT 624.0500 1119.3800 627.7500 1120.0000 ;
      RECT 620.0500 1119.3800 623.7500 1120.0000 ;
      RECT 616.0500 1119.3800 619.7500 1120.0000 ;
      RECT 612.0500 1119.3800 615.7500 1120.0000 ;
      RECT 608.0500 1119.3800 611.7500 1120.0000 ;
      RECT 604.0500 1119.3800 607.7500 1120.0000 ;
      RECT 600.0500 1119.3800 603.7500 1120.0000 ;
      RECT 596.0500 1119.3800 599.7500 1120.0000 ;
      RECT 592.0500 1119.3800 595.7500 1120.0000 ;
      RECT 588.0500 1119.3800 591.7500 1120.0000 ;
      RECT 584.0500 1119.3800 587.7500 1120.0000 ;
      RECT 580.0500 1119.3800 583.7500 1120.0000 ;
      RECT 576.0500 1119.3800 579.7500 1120.0000 ;
      RECT 572.0500 1119.3800 575.7500 1120.0000 ;
      RECT 568.0500 1119.3800 571.7500 1120.0000 ;
      RECT 564.0500 1119.3800 567.7500 1120.0000 ;
      RECT 560.0500 1119.3800 563.7500 1120.0000 ;
      RECT 556.0500 1119.3800 559.7500 1120.0000 ;
      RECT 552.0500 1119.3800 555.7500 1120.0000 ;
      RECT 548.0500 1119.3800 551.7500 1120.0000 ;
      RECT 544.0500 1119.3800 547.7500 1120.0000 ;
      RECT 540.0500 1119.3800 543.7500 1120.0000 ;
      RECT 536.0500 1119.3800 539.7500 1120.0000 ;
      RECT 532.0500 1119.3800 535.7500 1120.0000 ;
      RECT 528.0500 1119.3800 531.7500 1120.0000 ;
      RECT 524.0500 1119.3800 527.7500 1120.0000 ;
      RECT 520.0500 1119.3800 523.7500 1120.0000 ;
      RECT 516.0500 1119.3800 519.7500 1120.0000 ;
      RECT 512.0500 1119.3800 515.7500 1120.0000 ;
      RECT 508.0500 1119.3800 511.7500 1120.0000 ;
      RECT 504.0500 1119.3800 507.7500 1120.0000 ;
      RECT 500.0500 1119.3800 503.7500 1120.0000 ;
      RECT 496.0500 1119.3800 499.7500 1120.0000 ;
      RECT 492.0500 1119.3800 495.7500 1120.0000 ;
      RECT 488.0500 1119.3800 491.7500 1120.0000 ;
      RECT 484.0500 1119.3800 487.7500 1120.0000 ;
      RECT 480.0500 1119.3800 483.7500 1120.0000 ;
      RECT 476.0500 1119.3800 479.7500 1120.0000 ;
      RECT 472.0500 1119.3800 475.7500 1120.0000 ;
      RECT 468.0500 1119.3800 471.7500 1120.0000 ;
      RECT 464.0500 1119.3800 467.7500 1120.0000 ;
      RECT 460.0500 1119.3800 463.7500 1120.0000 ;
      RECT 456.0500 1119.3800 459.7500 1120.0000 ;
      RECT 452.0500 1119.3800 455.7500 1120.0000 ;
      RECT 448.0500 1119.3800 451.7500 1120.0000 ;
      RECT 444.0500 1119.3800 447.7500 1120.0000 ;
      RECT 440.0500 1119.3800 443.7500 1120.0000 ;
      RECT 436.0500 1119.3800 439.7500 1120.0000 ;
      RECT 432.0500 1119.3800 435.7500 1120.0000 ;
      RECT 428.0500 1119.3800 431.7500 1120.0000 ;
      RECT 424.0500 1119.3800 427.7500 1120.0000 ;
      RECT 420.0500 1119.3800 423.7500 1120.0000 ;
      RECT 416.0500 1119.3800 419.7500 1120.0000 ;
      RECT 412.0500 1119.3800 415.7500 1120.0000 ;
      RECT 408.0500 1119.3800 411.7500 1120.0000 ;
      RECT 404.0500 1119.3800 407.7500 1120.0000 ;
      RECT 400.0500 1119.3800 403.7500 1120.0000 ;
      RECT 396.0500 1119.3800 399.7500 1120.0000 ;
      RECT 0.0000 1119.3800 395.7500 1120.0000 ;
      RECT 0.0000 0.6200 1120.0000 1119.3800 ;
      RECT 926.2500 0.0000 1120.0000 0.6200 ;
      RECT 922.2500 0.0000 925.9500 0.6200 ;
      RECT 918.2500 0.0000 921.9500 0.6200 ;
      RECT 914.2500 0.0000 917.9500 0.6200 ;
      RECT 910.2500 0.0000 913.9500 0.6200 ;
      RECT 906.2500 0.0000 909.9500 0.6200 ;
      RECT 902.2500 0.0000 905.9500 0.6200 ;
      RECT 898.2500 0.0000 901.9500 0.6200 ;
      RECT 894.2500 0.0000 897.9500 0.6200 ;
      RECT 890.2500 0.0000 893.9500 0.6200 ;
      RECT 886.2500 0.0000 889.9500 0.6200 ;
      RECT 882.2500 0.0000 885.9500 0.6200 ;
      RECT 878.2500 0.0000 881.9500 0.6200 ;
      RECT 874.2500 0.0000 877.9500 0.6200 ;
      RECT 870.2500 0.0000 873.9500 0.6200 ;
      RECT 866.2500 0.0000 869.9500 0.6200 ;
      RECT 862.2500 0.0000 865.9500 0.6200 ;
      RECT 858.2500 0.0000 861.9500 0.6200 ;
      RECT 854.2500 0.0000 857.9500 0.6200 ;
      RECT 850.2500 0.0000 853.9500 0.6200 ;
      RECT 846.2500 0.0000 849.9500 0.6200 ;
      RECT 842.2500 0.0000 845.9500 0.6200 ;
      RECT 838.2500 0.0000 841.9500 0.6200 ;
      RECT 834.2500 0.0000 837.9500 0.6200 ;
      RECT 830.2500 0.0000 833.9500 0.6200 ;
      RECT 826.2500 0.0000 829.9500 0.6200 ;
      RECT 822.2500 0.0000 825.9500 0.6200 ;
      RECT 818.2500 0.0000 821.9500 0.6200 ;
      RECT 814.2500 0.0000 817.9500 0.6200 ;
      RECT 810.2500 0.0000 813.9500 0.6200 ;
      RECT 806.2500 0.0000 809.9500 0.6200 ;
      RECT 802.2500 0.0000 805.9500 0.6200 ;
      RECT 798.2500 0.0000 801.9500 0.6200 ;
      RECT 794.2500 0.0000 797.9500 0.6200 ;
      RECT 790.2500 0.0000 793.9500 0.6200 ;
      RECT 786.2500 0.0000 789.9500 0.6200 ;
      RECT 782.2500 0.0000 785.9500 0.6200 ;
      RECT 778.2500 0.0000 781.9500 0.6200 ;
      RECT 774.2500 0.0000 777.9500 0.6200 ;
      RECT 770.2500 0.0000 773.9500 0.6200 ;
      RECT 766.2500 0.0000 769.9500 0.6200 ;
      RECT 762.2500 0.0000 765.9500 0.6200 ;
      RECT 758.2500 0.0000 761.9500 0.6200 ;
      RECT 754.2500 0.0000 757.9500 0.6200 ;
      RECT 750.2500 0.0000 753.9500 0.6200 ;
      RECT 746.2500 0.0000 749.9500 0.6200 ;
      RECT 742.2500 0.0000 745.9500 0.6200 ;
      RECT 738.2500 0.0000 741.9500 0.6200 ;
      RECT 734.2500 0.0000 737.9500 0.6200 ;
      RECT 730.2500 0.0000 733.9500 0.6200 ;
      RECT 726.2500 0.0000 729.9500 0.6200 ;
      RECT 722.2500 0.0000 725.9500 0.6200 ;
      RECT 718.2500 0.0000 721.9500 0.6200 ;
      RECT 714.2500 0.0000 717.9500 0.6200 ;
      RECT 710.2500 0.0000 713.9500 0.6200 ;
      RECT 706.2500 0.0000 709.9500 0.6200 ;
      RECT 702.2500 0.0000 705.9500 0.6200 ;
      RECT 698.2500 0.0000 701.9500 0.6200 ;
      RECT 694.2500 0.0000 697.9500 0.6200 ;
      RECT 690.2500 0.0000 693.9500 0.6200 ;
      RECT 686.2500 0.0000 689.9500 0.6200 ;
      RECT 682.2500 0.0000 685.9500 0.6200 ;
      RECT 678.2500 0.0000 681.9500 0.6200 ;
      RECT 674.2500 0.0000 677.9500 0.6200 ;
      RECT 670.2500 0.0000 673.9500 0.6200 ;
      RECT 666.2500 0.0000 669.9500 0.6200 ;
      RECT 662.2500 0.0000 665.9500 0.6200 ;
      RECT 658.2500 0.0000 661.9500 0.6200 ;
      RECT 654.2500 0.0000 657.9500 0.6200 ;
      RECT 650.2500 0.0000 653.9500 0.6200 ;
      RECT 646.2500 0.0000 649.9500 0.6200 ;
      RECT 642.2500 0.0000 645.9500 0.6200 ;
      RECT 638.2500 0.0000 641.9500 0.6200 ;
      RECT 634.2500 0.0000 637.9500 0.6200 ;
      RECT 630.2500 0.0000 633.9500 0.6200 ;
      RECT 626.2500 0.0000 629.9500 0.6200 ;
      RECT 622.2500 0.0000 625.9500 0.6200 ;
      RECT 618.2500 0.0000 621.9500 0.6200 ;
      RECT 614.2500 0.0000 617.9500 0.6200 ;
      RECT 610.2500 0.0000 613.9500 0.6200 ;
      RECT 606.2500 0.0000 609.9500 0.6200 ;
      RECT 602.2500 0.0000 605.9500 0.6200 ;
      RECT 598.2500 0.0000 601.9500 0.6200 ;
      RECT 594.2500 0.0000 597.9500 0.6200 ;
      RECT 590.2500 0.0000 593.9500 0.6200 ;
      RECT 586.2500 0.0000 589.9500 0.6200 ;
      RECT 582.2500 0.0000 585.9500 0.6200 ;
      RECT 578.2500 0.0000 581.9500 0.6200 ;
      RECT 574.2500 0.0000 577.9500 0.6200 ;
      RECT 570.2500 0.0000 573.9500 0.6200 ;
      RECT 566.2500 0.0000 569.9500 0.6200 ;
      RECT 562.2500 0.0000 565.9500 0.6200 ;
      RECT 558.2500 0.0000 561.9500 0.6200 ;
      RECT 554.2500 0.0000 557.9500 0.6200 ;
      RECT 550.2500 0.0000 553.9500 0.6200 ;
      RECT 546.2500 0.0000 549.9500 0.6200 ;
      RECT 542.2500 0.0000 545.9500 0.6200 ;
      RECT 538.2500 0.0000 541.9500 0.6200 ;
      RECT 534.2500 0.0000 537.9500 0.6200 ;
      RECT 530.2500 0.0000 533.9500 0.6200 ;
      RECT 526.2500 0.0000 529.9500 0.6200 ;
      RECT 522.2500 0.0000 525.9500 0.6200 ;
      RECT 518.2500 0.0000 521.9500 0.6200 ;
      RECT 514.2500 0.0000 517.9500 0.6200 ;
      RECT 510.2500 0.0000 513.9500 0.6200 ;
      RECT 506.2500 0.0000 509.9500 0.6200 ;
      RECT 502.2500 0.0000 505.9500 0.6200 ;
      RECT 498.2500 0.0000 501.9500 0.6200 ;
      RECT 494.2500 0.0000 497.9500 0.6200 ;
      RECT 490.2500 0.0000 493.9500 0.6200 ;
      RECT 486.2500 0.0000 489.9500 0.6200 ;
      RECT 482.2500 0.0000 485.9500 0.6200 ;
      RECT 478.2500 0.0000 481.9500 0.6200 ;
      RECT 474.2500 0.0000 477.9500 0.6200 ;
      RECT 470.2500 0.0000 473.9500 0.6200 ;
      RECT 466.2500 0.0000 469.9500 0.6200 ;
      RECT 462.2500 0.0000 465.9500 0.6200 ;
      RECT 458.2500 0.0000 461.9500 0.6200 ;
      RECT 454.2500 0.0000 457.9500 0.6200 ;
      RECT 450.2500 0.0000 453.9500 0.6200 ;
      RECT 446.2500 0.0000 449.9500 0.6200 ;
      RECT 442.2500 0.0000 445.9500 0.6200 ;
      RECT 438.2500 0.0000 441.9500 0.6200 ;
      RECT 434.2500 0.0000 437.9500 0.6200 ;
      RECT 430.2500 0.0000 433.9500 0.6200 ;
      RECT 426.2500 0.0000 429.9500 0.6200 ;
      RECT 422.2500 0.0000 425.9500 0.6200 ;
      RECT 418.2500 0.0000 421.9500 0.6200 ;
      RECT 414.2500 0.0000 417.9500 0.6200 ;
      RECT 410.2500 0.0000 413.9500 0.6200 ;
      RECT 406.2500 0.0000 409.9500 0.6200 ;
      RECT 402.2500 0.0000 405.9500 0.6200 ;
      RECT 398.2500 0.0000 401.9500 0.6200 ;
      RECT 394.2500 0.0000 397.9500 0.6200 ;
      RECT 390.2500 0.0000 393.9500 0.6200 ;
      RECT 386.2500 0.0000 389.9500 0.6200 ;
      RECT 382.2500 0.0000 385.9500 0.6200 ;
      RECT 378.2500 0.0000 381.9500 0.6200 ;
      RECT 374.2500 0.0000 377.9500 0.6200 ;
      RECT 370.2500 0.0000 373.9500 0.6200 ;
      RECT 366.2500 0.0000 369.9500 0.6200 ;
      RECT 362.2500 0.0000 365.9500 0.6200 ;
      RECT 358.2500 0.0000 361.9500 0.6200 ;
      RECT 354.2500 0.0000 357.9500 0.6200 ;
      RECT 350.2500 0.0000 353.9500 0.6200 ;
      RECT 346.2500 0.0000 349.9500 0.6200 ;
      RECT 342.2500 0.0000 345.9500 0.6200 ;
      RECT 338.2500 0.0000 341.9500 0.6200 ;
      RECT 334.2500 0.0000 337.9500 0.6200 ;
      RECT 330.2500 0.0000 333.9500 0.6200 ;
      RECT 326.2500 0.0000 329.9500 0.6200 ;
      RECT 322.2500 0.0000 325.9500 0.6200 ;
      RECT 318.2500 0.0000 321.9500 0.6200 ;
      RECT 314.2500 0.0000 317.9500 0.6200 ;
      RECT 310.2500 0.0000 313.9500 0.6200 ;
      RECT 306.2500 0.0000 309.9500 0.6200 ;
      RECT 302.2500 0.0000 305.9500 0.6200 ;
      RECT 298.2500 0.0000 301.9500 0.6200 ;
      RECT 294.2500 0.0000 297.9500 0.6200 ;
      RECT 290.2500 0.0000 293.9500 0.6200 ;
      RECT 286.2500 0.0000 289.9500 0.6200 ;
      RECT 282.2500 0.0000 285.9500 0.6200 ;
      RECT 278.2500 0.0000 281.9500 0.6200 ;
      RECT 274.2500 0.0000 277.9500 0.6200 ;
      RECT 270.2500 0.0000 273.9500 0.6200 ;
      RECT 266.2500 0.0000 269.9500 0.6200 ;
      RECT 262.2500 0.0000 265.9500 0.6200 ;
      RECT 258.2500 0.0000 261.9500 0.6200 ;
      RECT 254.2500 0.0000 257.9500 0.6200 ;
      RECT 250.2500 0.0000 253.9500 0.6200 ;
      RECT 246.2500 0.0000 249.9500 0.6200 ;
      RECT 242.2500 0.0000 245.9500 0.6200 ;
      RECT 238.2500 0.0000 241.9500 0.6200 ;
      RECT 234.2500 0.0000 237.9500 0.6200 ;
      RECT 230.2500 0.0000 233.9500 0.6200 ;
      RECT 226.2500 0.0000 229.9500 0.6200 ;
      RECT 222.2500 0.0000 225.9500 0.6200 ;
      RECT 218.2500 0.0000 221.9500 0.6200 ;
      RECT 214.2500 0.0000 217.9500 0.6200 ;
      RECT 210.2500 0.0000 213.9500 0.6200 ;
      RECT 206.2500 0.0000 209.9500 0.6200 ;
      RECT 202.2500 0.0000 205.9500 0.6200 ;
      RECT 198.2500 0.0000 201.9500 0.6200 ;
      RECT 194.2500 0.0000 197.9500 0.6200 ;
      RECT 0.0000 0.0000 193.9500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 1120.0000 1120.0000 ;
    LAYER M4 ;
      RECT 0.0000 1118.4000 1120.0000 1120.0000 ;
      RECT 0.0000 1110.1300 1114.0000 1118.4000 ;
      RECT 8.5000 1107.1300 1111.5000 1110.1300 ;
      RECT 0.0000 1107.1300 5.5000 1110.1300 ;
      RECT 1117.0000 1105.1300 1120.0000 1118.4000 ;
      RECT 0.0000 1103.0350 1114.0000 1107.1300 ;
      RECT 1118.5000 1102.1300 1120.0000 1105.1300 ;
      RECT 8.5000 1100.0350 1111.5000 1103.0350 ;
      RECT 0.0000 1100.0350 5.5000 1103.0350 ;
      RECT 1117.0000 1098.0350 1120.0000 1102.1300 ;
      RECT 0.0000 1095.9400 1114.0000 1100.0350 ;
      RECT 1118.5000 1095.0350 1120.0000 1098.0350 ;
      RECT 8.5000 1092.9400 1111.5000 1095.9400 ;
      RECT 0.0000 1092.9400 5.5000 1095.9400 ;
      RECT 1117.0000 1090.9400 1120.0000 1095.0350 ;
      RECT 0.0000 1088.8450 1114.0000 1092.9400 ;
      RECT 1118.5000 1087.9400 1120.0000 1090.9400 ;
      RECT 8.5000 1085.8450 1111.5000 1088.8450 ;
      RECT 0.0000 1085.8450 5.5000 1088.8450 ;
      RECT 1117.0000 1083.8450 1120.0000 1087.9400 ;
      RECT 0.0000 1081.7500 1114.0000 1085.8450 ;
      RECT 1118.5000 1080.8450 1120.0000 1083.8450 ;
      RECT 8.5000 1078.7500 1111.5000 1081.7500 ;
      RECT 0.0000 1078.7500 5.5000 1081.7500 ;
      RECT 1117.0000 1076.7500 1120.0000 1080.8450 ;
      RECT 0.0000 1074.6550 1114.0000 1078.7500 ;
      RECT 1118.5000 1073.7500 1120.0000 1076.7500 ;
      RECT 8.5000 1071.6550 1111.5000 1074.6550 ;
      RECT 0.0000 1071.6550 5.5000 1074.6550 ;
      RECT 1117.0000 1069.6550 1120.0000 1073.7500 ;
      RECT 0.0000 1067.5600 1114.0000 1071.6550 ;
      RECT 1118.5000 1066.6550 1120.0000 1069.6550 ;
      RECT 8.5000 1064.5600 1111.5000 1067.5600 ;
      RECT 0.0000 1064.5600 5.5000 1067.5600 ;
      RECT 1117.0000 1062.5600 1120.0000 1066.6550 ;
      RECT 0.0000 1060.4650 1114.0000 1064.5600 ;
      RECT 1118.5000 1059.5600 1120.0000 1062.5600 ;
      RECT 8.5000 1057.4650 1111.5000 1060.4650 ;
      RECT 0.0000 1057.4650 5.5000 1060.4650 ;
      RECT 1117.0000 1055.4650 1120.0000 1059.5600 ;
      RECT 0.0000 1053.3700 1114.0000 1057.4650 ;
      RECT 1118.5000 1052.4650 1120.0000 1055.4650 ;
      RECT 8.5000 1050.3700 1111.5000 1053.3700 ;
      RECT 0.0000 1050.3700 5.5000 1053.3700 ;
      RECT 1117.0000 1048.3700 1120.0000 1052.4650 ;
      RECT 0.0000 1046.2750 1114.0000 1050.3700 ;
      RECT 1118.5000 1045.3700 1120.0000 1048.3700 ;
      RECT 8.5000 1043.2750 1111.5000 1046.2750 ;
      RECT 0.0000 1043.2750 5.5000 1046.2750 ;
      RECT 1117.0000 1041.2750 1120.0000 1045.3700 ;
      RECT 0.0000 1039.1800 1114.0000 1043.2750 ;
      RECT 1118.5000 1038.2750 1120.0000 1041.2750 ;
      RECT 8.5000 1036.1800 1111.5000 1039.1800 ;
      RECT 0.0000 1036.1800 5.5000 1039.1800 ;
      RECT 1117.0000 1034.1800 1120.0000 1038.2750 ;
      RECT 0.0000 1032.0850 1114.0000 1036.1800 ;
      RECT 1118.5000 1031.1800 1120.0000 1034.1800 ;
      RECT 8.5000 1029.0850 1111.5000 1032.0850 ;
      RECT 0.0000 1029.0850 5.5000 1032.0850 ;
      RECT 1117.0000 1027.0850 1120.0000 1031.1800 ;
      RECT 0.0000 1024.9900 1114.0000 1029.0850 ;
      RECT 1118.5000 1024.0850 1120.0000 1027.0850 ;
      RECT 8.5000 1021.9900 1111.5000 1024.9900 ;
      RECT 0.0000 1021.9900 5.5000 1024.9900 ;
      RECT 1117.0000 1019.9900 1120.0000 1024.0850 ;
      RECT 0.0000 1017.8950 1114.0000 1021.9900 ;
      RECT 1118.5000 1016.9900 1120.0000 1019.9900 ;
      RECT 8.5000 1014.8950 1111.5000 1017.8950 ;
      RECT 0.0000 1014.8950 5.5000 1017.8950 ;
      RECT 1117.0000 1012.8950 1120.0000 1016.9900 ;
      RECT 0.0000 1010.8000 1114.0000 1014.8950 ;
      RECT 1118.5000 1009.8950 1120.0000 1012.8950 ;
      RECT 1114.5000 1007.8000 1120.0000 1009.8950 ;
      RECT 8.5000 1007.8000 1111.5000 1010.8000 ;
      RECT 0.0000 1007.8000 5.5000 1010.8000 ;
      RECT 0.0000 1005.8000 1120.0000 1007.8000 ;
      RECT 4.5000 1003.9250 1115.5000 1005.8000 ;
      RECT 4.5000 1003.7050 1114.5550 1003.9250 ;
      RECT 1115.2850 1003.2750 1115.5000 1003.9250 ;
      RECT 1114.5000 1003.2750 1114.5550 1003.7050 ;
      RECT 1118.5000 1002.8000 1120.0000 1005.8000 ;
      RECT 1114.5000 1002.8000 1115.5000 1003.2750 ;
      RECT 4.5000 1002.8000 5.5000 1003.7050 ;
      RECT 0.0000 1002.8000 1.5000 1005.8000 ;
      RECT 1114.5000 1000.7050 1120.0000 1002.8000 ;
      RECT 8.5000 1000.7050 1111.5000 1003.7050 ;
      RECT 0.0000 1000.7050 5.5000 1002.8000 ;
      RECT 0.0000 998.7050 1120.0000 1000.7050 ;
      RECT 4.5000 996.7250 1115.5000 998.7050 ;
      RECT 4.5000 996.6100 1114.5550 996.7250 ;
      RECT 1115.2850 996.0750 1115.5000 996.7250 ;
      RECT 1114.5000 996.0750 1114.5550 996.6100 ;
      RECT 1118.5000 995.7050 1120.0000 998.7050 ;
      RECT 1114.5000 995.7050 1115.5000 996.0750 ;
      RECT 4.5000 995.7050 5.5000 996.6100 ;
      RECT 0.0000 995.7050 1.5000 998.7050 ;
      RECT 1114.5000 993.6100 1120.0000 995.7050 ;
      RECT 8.5000 993.6100 1111.5000 996.6100 ;
      RECT 0.0000 993.6100 5.5000 995.7050 ;
      RECT 0.0000 991.6100 1120.0000 993.6100 ;
      RECT 4.5000 989.5150 1115.5000 991.6100 ;
      RECT 1118.5000 988.6100 1120.0000 991.6100 ;
      RECT 1114.5000 988.6100 1115.5000 989.5150 ;
      RECT 4.5000 988.6100 5.5000 989.5150 ;
      RECT 0.0000 988.6100 1.5000 991.6100 ;
      RECT 1114.5000 986.5150 1120.0000 988.6100 ;
      RECT 8.5000 986.5150 1111.5000 989.5150 ;
      RECT 0.0000 986.5150 5.5000 988.6100 ;
      RECT 0.0000 984.5150 1120.0000 986.5150 ;
      RECT 4.5000 982.4200 1115.5000 984.5150 ;
      RECT 1118.5000 981.5150 1120.0000 984.5150 ;
      RECT 1114.5000 981.5150 1115.5000 982.4200 ;
      RECT 4.5000 981.5150 5.5000 982.4200 ;
      RECT 0.0000 981.5150 1.5000 984.5150 ;
      RECT 1114.5000 979.4200 1120.0000 981.5150 ;
      RECT 8.5000 979.4200 1111.5000 982.4200 ;
      RECT 0.0000 979.4200 5.5000 981.5150 ;
      RECT 0.0000 977.4200 1120.0000 979.4200 ;
      RECT 4.5000 975.3250 1115.5000 977.4200 ;
      RECT 1118.5000 974.4200 1120.0000 977.4200 ;
      RECT 1114.5000 974.4200 1115.5000 975.3250 ;
      RECT 4.5000 974.4200 5.5000 975.3250 ;
      RECT 0.0000 974.4200 1.5000 977.4200 ;
      RECT 1114.5000 972.3250 1120.0000 974.4200 ;
      RECT 8.5000 972.3250 1111.5000 975.3250 ;
      RECT 0.0000 972.3250 5.5000 974.4200 ;
      RECT 0.0000 970.3250 1120.0000 972.3250 ;
      RECT 4.5000 968.2300 1115.5000 970.3250 ;
      RECT 1118.5000 967.3250 1120.0000 970.3250 ;
      RECT 1114.5000 967.3250 1115.5000 968.2300 ;
      RECT 4.5000 967.3250 5.5000 968.2300 ;
      RECT 0.0000 967.3250 1.5000 970.3250 ;
      RECT 1114.5000 965.2300 1120.0000 967.3250 ;
      RECT 8.5000 965.2300 1111.5000 968.2300 ;
      RECT 0.0000 965.2300 5.5000 967.3250 ;
      RECT 0.0000 963.2300 1120.0000 965.2300 ;
      RECT 4.5000 961.1350 1115.5000 963.2300 ;
      RECT 1118.5000 960.2300 1120.0000 963.2300 ;
      RECT 1114.5000 960.2300 1115.5000 961.1350 ;
      RECT 4.5000 960.2300 5.5000 961.1350 ;
      RECT 0.0000 960.2300 1.5000 963.2300 ;
      RECT 1114.5000 958.1350 1120.0000 960.2300 ;
      RECT 8.5000 958.1350 1111.5000 961.1350 ;
      RECT 0.0000 958.1350 5.5000 960.2300 ;
      RECT 0.0000 956.1350 1120.0000 958.1350 ;
      RECT 4.5000 954.0400 1115.5000 956.1350 ;
      RECT 1118.5000 953.1350 1120.0000 956.1350 ;
      RECT 1114.5000 953.1350 1115.5000 954.0400 ;
      RECT 4.5000 953.1350 5.5000 954.0400 ;
      RECT 0.0000 953.1350 1.5000 956.1350 ;
      RECT 1114.5000 951.0400 1120.0000 953.1350 ;
      RECT 8.5000 951.0400 1111.5000 954.0400 ;
      RECT 0.0000 951.0400 5.5000 953.1350 ;
      RECT 0.0000 949.0400 1120.0000 951.0400 ;
      RECT 4.5000 946.9450 1115.5000 949.0400 ;
      RECT 1118.5000 946.0400 1120.0000 949.0400 ;
      RECT 1114.5000 946.0400 1115.5000 946.9450 ;
      RECT 4.5000 946.0400 5.5000 946.9450 ;
      RECT 0.0000 946.0400 1.5000 949.0400 ;
      RECT 1114.5000 943.9450 1120.0000 946.0400 ;
      RECT 8.5000 943.9450 1111.5000 946.9450 ;
      RECT 0.0000 943.9450 5.5000 946.0400 ;
      RECT 0.0000 941.9450 1120.0000 943.9450 ;
      RECT 4.5000 939.8500 1115.5000 941.9450 ;
      RECT 1118.5000 938.9450 1120.0000 941.9450 ;
      RECT 1114.5000 938.9450 1115.5000 939.8500 ;
      RECT 4.5000 938.9450 5.5000 939.8500 ;
      RECT 0.0000 938.9450 1.5000 941.9450 ;
      RECT 1114.5000 936.8500 1120.0000 938.9450 ;
      RECT 8.5000 936.8500 1111.5000 939.8500 ;
      RECT 0.0000 936.8500 5.5000 938.9450 ;
      RECT 0.0000 934.8500 1120.0000 936.8500 ;
      RECT 4.5000 932.7550 1115.5000 934.8500 ;
      RECT 1118.5000 931.8500 1120.0000 934.8500 ;
      RECT 1114.5000 931.8500 1115.5000 932.7550 ;
      RECT 4.5000 931.8500 5.5000 932.7550 ;
      RECT 0.0000 931.8500 1.5000 934.8500 ;
      RECT 1114.5000 929.7550 1120.0000 931.8500 ;
      RECT 8.5000 929.7550 1111.5000 932.7550 ;
      RECT 0.0000 929.7550 5.5000 931.8500 ;
      RECT 0.0000 927.7550 1120.0000 929.7550 ;
      RECT 4.5000 925.6600 1115.5000 927.7550 ;
      RECT 1118.5000 924.7550 1120.0000 927.7550 ;
      RECT 1114.5000 924.7550 1115.5000 925.6600 ;
      RECT 4.5000 924.7550 5.5000 925.6600 ;
      RECT 0.0000 924.7550 1.5000 927.7550 ;
      RECT 1114.5000 922.6600 1120.0000 924.7550 ;
      RECT 8.5000 922.6600 1111.5000 925.6600 ;
      RECT 0.0000 922.6600 5.5000 924.7550 ;
      RECT 0.0000 920.6600 1120.0000 922.6600 ;
      RECT 4.5000 918.5650 1115.5000 920.6600 ;
      RECT 1118.5000 917.6600 1120.0000 920.6600 ;
      RECT 1114.5000 917.6600 1115.5000 918.5650 ;
      RECT 4.5000 917.6600 5.5000 918.5650 ;
      RECT 0.0000 917.6600 1.5000 920.6600 ;
      RECT 1114.5000 915.5650 1120.0000 917.6600 ;
      RECT 8.5000 915.5650 1111.5000 918.5650 ;
      RECT 0.0000 915.5650 5.5000 917.6600 ;
      RECT 0.0000 913.5650 1120.0000 915.5650 ;
      RECT 4.5000 911.4700 1115.5000 913.5650 ;
      RECT 1118.5000 910.5650 1120.0000 913.5650 ;
      RECT 1114.5000 910.5650 1115.5000 911.4700 ;
      RECT 4.5000 910.5650 5.5000 911.4700 ;
      RECT 0.0000 910.5650 1.5000 913.5650 ;
      RECT 1114.5000 908.4700 1120.0000 910.5650 ;
      RECT 8.5000 908.4700 1111.5000 911.4700 ;
      RECT 0.0000 908.4700 5.5000 910.5650 ;
      RECT 0.0000 906.4700 1120.0000 908.4700 ;
      RECT 4.5000 904.3750 1115.5000 906.4700 ;
      RECT 1118.5000 903.4700 1120.0000 906.4700 ;
      RECT 1114.5000 903.4700 1115.5000 904.3750 ;
      RECT 4.5000 903.4700 5.5000 904.3750 ;
      RECT 0.0000 903.4700 1.5000 906.4700 ;
      RECT 1114.5000 901.3750 1120.0000 903.4700 ;
      RECT 8.5000 901.3750 1111.5000 904.3750 ;
      RECT 0.0000 901.3750 5.5000 903.4700 ;
      RECT 0.0000 899.3750 1120.0000 901.3750 ;
      RECT 4.5000 897.2800 1115.5000 899.3750 ;
      RECT 1118.5000 896.3750 1120.0000 899.3750 ;
      RECT 1114.5000 896.3750 1115.5000 897.2800 ;
      RECT 4.5000 896.3750 5.5000 897.2800 ;
      RECT 0.0000 896.3750 1.5000 899.3750 ;
      RECT 1114.5000 894.2800 1120.0000 896.3750 ;
      RECT 8.5000 894.2800 1111.5000 897.2800 ;
      RECT 0.0000 894.2800 5.5000 896.3750 ;
      RECT 0.0000 892.2800 1120.0000 894.2800 ;
      RECT 4.5000 890.1850 1115.5000 892.2800 ;
      RECT 1118.5000 889.2800 1120.0000 892.2800 ;
      RECT 1114.5000 889.2800 1115.5000 890.1850 ;
      RECT 4.5000 889.2800 5.5000 890.1850 ;
      RECT 0.0000 889.2800 1.5000 892.2800 ;
      RECT 1114.5000 887.1850 1120.0000 889.2800 ;
      RECT 8.5000 887.1850 1111.5000 890.1850 ;
      RECT 0.0000 887.1850 5.5000 889.2800 ;
      RECT 0.0000 885.1850 1120.0000 887.1850 ;
      RECT 4.5000 883.0900 1115.5000 885.1850 ;
      RECT 1118.5000 882.1850 1120.0000 885.1850 ;
      RECT 1114.5000 882.1850 1115.5000 883.0900 ;
      RECT 4.5000 882.1850 5.5000 883.0900 ;
      RECT 0.0000 882.1850 1.5000 885.1850 ;
      RECT 1114.5000 880.0900 1120.0000 882.1850 ;
      RECT 8.5000 880.0900 1111.5000 883.0900 ;
      RECT 0.0000 880.0900 5.5000 882.1850 ;
      RECT 0.0000 878.0900 1120.0000 880.0900 ;
      RECT 4.5000 875.9950 1115.5000 878.0900 ;
      RECT 1118.5000 875.0900 1120.0000 878.0900 ;
      RECT 1114.5000 875.0900 1115.5000 875.9950 ;
      RECT 4.5000 875.0900 5.5000 875.9950 ;
      RECT 0.0000 875.0900 1.5000 878.0900 ;
      RECT 1114.5000 872.9950 1120.0000 875.0900 ;
      RECT 8.5000 872.9950 1111.5000 875.9950 ;
      RECT 0.0000 872.9950 5.5000 875.0900 ;
      RECT 0.0000 870.9950 1120.0000 872.9950 ;
      RECT 4.5000 868.9000 1115.5000 870.9950 ;
      RECT 1118.5000 867.9950 1120.0000 870.9950 ;
      RECT 1114.5000 867.9950 1115.5000 868.9000 ;
      RECT 4.5000 867.9950 5.5000 868.9000 ;
      RECT 0.0000 867.9950 1.5000 870.9950 ;
      RECT 1114.5000 865.9000 1120.0000 867.9950 ;
      RECT 8.5000 865.9000 1111.5000 868.9000 ;
      RECT 0.0000 865.9000 5.5000 867.9950 ;
      RECT 0.0000 863.9000 1120.0000 865.9000 ;
      RECT 4.5000 863.5250 1115.5000 863.9000 ;
      RECT 1115.2850 862.8750 1115.5000 863.5250 ;
      RECT 4.5000 862.8750 1114.5550 863.5250 ;
      RECT 4.5000 861.8050 1115.5000 862.8750 ;
      RECT 1118.5000 860.9000 1120.0000 863.9000 ;
      RECT 1114.5000 860.9000 1115.5000 861.8050 ;
      RECT 4.5000 860.9000 5.5000 861.8050 ;
      RECT 0.0000 860.9000 1.5000 863.9000 ;
      RECT 1114.5000 858.8050 1120.0000 860.9000 ;
      RECT 8.5000 858.8050 1111.5000 861.8050 ;
      RECT 0.0000 858.8050 5.5000 860.9000 ;
      RECT 0.0000 856.8050 1120.0000 858.8050 ;
      RECT 4.5000 856.3250 1115.5000 856.8050 ;
      RECT 1115.2850 855.6750 1115.5000 856.3250 ;
      RECT 4.5000 855.6750 1114.5550 856.3250 ;
      RECT 4.5000 854.7100 1115.5000 855.6750 ;
      RECT 1118.5000 853.8050 1120.0000 856.8050 ;
      RECT 1114.5000 853.8050 1115.5000 854.7100 ;
      RECT 4.5000 853.8050 5.5000 854.7100 ;
      RECT 0.0000 853.8050 1.5000 856.8050 ;
      RECT 1114.5000 851.7100 1120.0000 853.8050 ;
      RECT 8.5000 851.7100 1111.5000 854.7100 ;
      RECT 0.0000 851.7100 5.5000 853.8050 ;
      RECT 0.0000 849.7100 1120.0000 851.7100 ;
      RECT 4.5000 849.1250 1115.5000 849.7100 ;
      RECT 1115.2850 848.4750 1115.5000 849.1250 ;
      RECT 4.5000 848.4750 1114.5550 849.1250 ;
      RECT 4.5000 847.6150 1115.5000 848.4750 ;
      RECT 1118.5000 846.7100 1120.0000 849.7100 ;
      RECT 1114.5000 846.7100 1115.5000 847.6150 ;
      RECT 4.5000 846.7100 5.5000 847.6150 ;
      RECT 0.0000 846.7100 1.5000 849.7100 ;
      RECT 1114.5000 844.6150 1120.0000 846.7100 ;
      RECT 8.5000 844.6150 1111.5000 847.6150 ;
      RECT 0.0000 844.6150 5.5000 846.7100 ;
      RECT 0.0000 842.6150 1120.0000 844.6150 ;
      RECT 4.5000 841.9250 1115.5000 842.6150 ;
      RECT 1115.2850 841.2750 1115.5000 841.9250 ;
      RECT 4.5000 841.2750 1114.5550 841.9250 ;
      RECT 4.5000 840.5200 1115.5000 841.2750 ;
      RECT 1118.5000 839.6150 1120.0000 842.6150 ;
      RECT 1114.5000 839.6150 1115.5000 840.5200 ;
      RECT 4.5000 839.6150 5.5000 840.5200 ;
      RECT 0.0000 839.6150 1.5000 842.6150 ;
      RECT 1114.5000 837.5200 1120.0000 839.6150 ;
      RECT 8.5000 837.5200 1111.5000 840.5200 ;
      RECT 0.0000 837.5200 5.5000 839.6150 ;
      RECT 0.0000 835.5200 1120.0000 837.5200 ;
      RECT 4.5000 834.7250 1115.5000 835.5200 ;
      RECT 1115.2850 834.0750 1115.5000 834.7250 ;
      RECT 4.5000 834.0750 1114.5550 834.7250 ;
      RECT 4.5000 833.4250 1115.5000 834.0750 ;
      RECT 1118.5000 832.5200 1120.0000 835.5200 ;
      RECT 1114.5000 832.5200 1115.5000 833.4250 ;
      RECT 4.5000 832.5200 5.5000 833.4250 ;
      RECT 0.0000 832.5200 1.5000 835.5200 ;
      RECT 1114.5000 830.4250 1120.0000 832.5200 ;
      RECT 8.5000 830.4250 1111.5000 833.4250 ;
      RECT 0.0000 830.4250 5.5000 832.5200 ;
      RECT 0.0000 828.4250 1120.0000 830.4250 ;
      RECT 4.5000 827.5250 1115.5000 828.4250 ;
      RECT 1115.2850 826.8750 1115.5000 827.5250 ;
      RECT 4.5000 826.8750 1114.5550 827.5250 ;
      RECT 4.5000 826.3300 1115.5000 826.8750 ;
      RECT 1118.5000 825.4250 1120.0000 828.4250 ;
      RECT 1114.5000 825.4250 1115.5000 826.3300 ;
      RECT 4.5000 825.4250 5.5000 826.3300 ;
      RECT 0.0000 825.4250 1.5000 828.4250 ;
      RECT 1114.5000 823.3300 1120.0000 825.4250 ;
      RECT 8.5000 823.3300 1111.5000 826.3300 ;
      RECT 0.0000 823.3300 5.5000 825.4250 ;
      RECT 0.0000 821.3300 1120.0000 823.3300 ;
      RECT 4.5000 820.3250 1115.5000 821.3300 ;
      RECT 1115.2850 819.6750 1115.5000 820.3250 ;
      RECT 4.5000 819.6750 1114.5550 820.3250 ;
      RECT 4.5000 819.2350 1115.5000 819.6750 ;
      RECT 1118.5000 818.3300 1120.0000 821.3300 ;
      RECT 1114.5000 818.3300 1115.5000 819.2350 ;
      RECT 4.5000 818.3300 5.5000 819.2350 ;
      RECT 0.0000 818.3300 1.5000 821.3300 ;
      RECT 1114.5000 816.2350 1120.0000 818.3300 ;
      RECT 8.5000 816.2350 1111.5000 819.2350 ;
      RECT 0.0000 816.2350 5.5000 818.3300 ;
      RECT 0.0000 814.2350 1120.0000 816.2350 ;
      RECT 4.5000 813.1250 1115.5000 814.2350 ;
      RECT 1115.2850 812.4750 1115.5000 813.1250 ;
      RECT 4.5000 812.4750 1114.5550 813.1250 ;
      RECT 4.5000 812.1400 1115.5000 812.4750 ;
      RECT 1118.5000 811.2350 1120.0000 814.2350 ;
      RECT 1114.5000 811.2350 1115.5000 812.1400 ;
      RECT 4.5000 811.2350 5.5000 812.1400 ;
      RECT 0.0000 811.2350 1.5000 814.2350 ;
      RECT 1114.5000 809.1400 1120.0000 811.2350 ;
      RECT 8.5000 809.1400 1111.5000 812.1400 ;
      RECT 0.0000 809.1400 5.5000 811.2350 ;
      RECT 0.0000 807.1400 1120.0000 809.1400 ;
      RECT 4.5000 805.9250 1115.5000 807.1400 ;
      RECT 1115.2850 805.2750 1115.5000 805.9250 ;
      RECT 4.5000 805.2750 1114.5550 805.9250 ;
      RECT 4.5000 805.0450 1115.5000 805.2750 ;
      RECT 1118.5000 804.1400 1120.0000 807.1400 ;
      RECT 1114.5000 804.1400 1115.5000 805.0450 ;
      RECT 4.5000 804.1400 5.5000 805.0450 ;
      RECT 0.0000 804.1400 1.5000 807.1400 ;
      RECT 1114.5000 802.0450 1120.0000 804.1400 ;
      RECT 8.5000 802.0450 1111.5000 805.0450 ;
      RECT 0.0000 802.0450 5.5000 804.1400 ;
      RECT 0.0000 800.0450 1120.0000 802.0450 ;
      RECT 4.5000 798.7250 1115.5000 800.0450 ;
      RECT 1115.2850 798.0750 1115.5000 798.7250 ;
      RECT 4.5000 798.0750 1114.5550 798.7250 ;
      RECT 4.5000 797.9500 1115.5000 798.0750 ;
      RECT 1118.5000 797.0450 1120.0000 800.0450 ;
      RECT 1114.5000 797.0450 1115.5000 797.9500 ;
      RECT 4.5000 797.0450 5.5000 797.9500 ;
      RECT 0.0000 797.0450 1.5000 800.0450 ;
      RECT 1114.5000 794.9500 1120.0000 797.0450 ;
      RECT 8.5000 794.9500 1111.5000 797.9500 ;
      RECT 0.0000 794.9500 5.5000 797.0450 ;
      RECT 0.0000 792.9500 1120.0000 794.9500 ;
      RECT 4.5000 791.5250 1115.5000 792.9500 ;
      RECT 1115.2850 790.8750 1115.5000 791.5250 ;
      RECT 4.5000 790.8750 1114.5550 791.5250 ;
      RECT 4.5000 790.8550 1115.5000 790.8750 ;
      RECT 1118.5000 789.9500 1120.0000 792.9500 ;
      RECT 1114.5000 789.9500 1115.5000 790.8550 ;
      RECT 4.5000 789.9500 5.5000 790.8550 ;
      RECT 0.0000 789.9500 1.5000 792.9500 ;
      RECT 1114.5000 787.8550 1120.0000 789.9500 ;
      RECT 8.5000 787.8550 1111.5000 790.8550 ;
      RECT 0.0000 787.8550 5.5000 789.9500 ;
      RECT 0.0000 785.8550 1120.0000 787.8550 ;
      RECT 0.0000 783.7600 1114.0000 785.8550 ;
      RECT 1118.5000 782.8550 1120.0000 785.8550 ;
      RECT 8.5000 780.7600 1111.5000 783.7600 ;
      RECT 0.0000 780.7600 5.5000 783.7600 ;
      RECT 1117.0000 778.7600 1120.0000 782.8550 ;
      RECT 0.0000 776.6650 1114.0000 780.7600 ;
      RECT 1118.5000 775.7600 1120.0000 778.7600 ;
      RECT 8.5000 773.6650 1111.5000 776.6650 ;
      RECT 0.0000 773.6650 5.5000 776.6650 ;
      RECT 1117.0000 771.6650 1120.0000 775.7600 ;
      RECT 0.0000 769.5700 1114.0000 773.6650 ;
      RECT 1118.5000 768.6650 1120.0000 771.6650 ;
      RECT 8.5000 766.5700 1111.5000 769.5700 ;
      RECT 0.0000 766.5700 5.5000 769.5700 ;
      RECT 1117.0000 764.5700 1120.0000 768.6650 ;
      RECT 0.0000 762.4750 1114.0000 766.5700 ;
      RECT 1118.5000 761.5700 1120.0000 764.5700 ;
      RECT 8.5000 759.4750 1111.5000 762.4750 ;
      RECT 0.0000 759.4750 5.5000 762.4750 ;
      RECT 1117.0000 757.4750 1120.0000 761.5700 ;
      RECT 0.0000 755.3800 1114.0000 759.4750 ;
      RECT 1118.5000 754.4750 1120.0000 757.4750 ;
      RECT 8.5000 752.3800 1111.5000 755.3800 ;
      RECT 0.0000 752.3800 5.5000 755.3800 ;
      RECT 1117.0000 750.3800 1120.0000 754.4750 ;
      RECT 0.0000 748.2850 1114.0000 752.3800 ;
      RECT 1118.5000 747.3800 1120.0000 750.3800 ;
      RECT 8.5000 745.2850 1111.5000 748.2850 ;
      RECT 0.0000 745.2850 5.5000 748.2850 ;
      RECT 1117.0000 743.2850 1120.0000 747.3800 ;
      RECT 0.0000 741.1900 1114.0000 745.2850 ;
      RECT 1118.5000 740.2850 1120.0000 743.2850 ;
      RECT 8.5000 738.1900 1111.5000 741.1900 ;
      RECT 0.0000 738.1900 5.5000 741.1900 ;
      RECT 1117.0000 736.1900 1120.0000 740.2850 ;
      RECT 0.0000 734.0950 1114.0000 738.1900 ;
      RECT 1118.5000 733.1900 1120.0000 736.1900 ;
      RECT 8.5000 731.0950 1111.5000 734.0950 ;
      RECT 0.0000 731.0950 5.5000 734.0950 ;
      RECT 1117.0000 729.0950 1120.0000 733.1900 ;
      RECT 0.0000 727.0000 1114.0000 731.0950 ;
      RECT 8.5000 726.5000 1111.5000 727.0000 ;
      RECT 1118.5000 726.0950 1120.0000 729.0950 ;
      RECT 1076.5000 724.0000 1111.5000 726.5000 ;
      RECT 396.5000 724.0000 1073.5000 726.5000 ;
      RECT 8.5000 724.0000 393.5000 726.5000 ;
      RECT 0.0000 724.0000 5.5000 727.0000 ;
      RECT 0.0000 723.5000 1114.0000 724.0000 ;
      RECT 412.6500 722.5000 1114.0000 723.5000 ;
      RECT 1117.0000 722.0000 1120.0000 726.0950 ;
      RECT 412.6500 720.5000 1113.6000 722.5000 ;
      RECT 0.0000 720.5000 409.6500 723.5000 ;
      RECT 0.0000 719.9050 1113.6000 720.5000 ;
      RECT 1118.5000 719.0000 1120.0000 722.0000 ;
      RECT 1114.5000 716.9050 1120.0000 719.0000 ;
      RECT 1076.5000 716.9050 1111.5000 719.9050 ;
      RECT 396.5000 716.9050 1073.5000 719.9050 ;
      RECT 8.5000 716.9050 393.5000 719.9050 ;
      RECT 0.0000 716.9050 5.5000 719.9050 ;
      RECT 0.0000 715.5000 1120.0000 716.9050 ;
      RECT 1116.6000 714.9050 1120.0000 715.5000 ;
      RECT 0.0000 712.8100 1113.6000 715.5000 ;
      RECT 1118.5000 711.9050 1120.0000 714.9050 ;
      RECT 396.5000 710.5000 1073.5000 712.8100 ;
      RECT 396.5000 710.3100 1057.5000 710.5000 ;
      RECT 1114.5000 709.8100 1120.0000 711.9050 ;
      RECT 1076.5000 709.8100 1111.5000 712.8100 ;
      RECT 1060.5000 709.8100 1073.5000 710.5000 ;
      RECT 396.5000 709.8100 409.6500 710.3100 ;
      RECT 8.5000 709.8100 393.5000 712.8100 ;
      RECT 0.0000 709.8100 5.5000 712.8100 ;
      RECT 1060.5000 708.3000 1120.0000 709.8100 ;
      RECT 1116.6000 707.8100 1120.0000 708.3000 ;
      RECT 412.6500 707.6650 1057.5000 710.3100 ;
      RECT 0.0000 707.6650 409.6500 709.8100 ;
      RECT 1060.5000 707.5000 1113.6000 708.3000 ;
      RECT 0.0000 707.5000 1057.5000 707.6650 ;
      RECT 0.0000 705.7150 1113.6000 707.5000 ;
      RECT 1118.5000 704.8100 1120.0000 707.8100 ;
      RECT 1114.5000 702.7150 1120.0000 704.8100 ;
      RECT 1076.5000 702.7150 1111.5000 705.7150 ;
      RECT 1060.5000 702.7150 1073.5000 705.7150 ;
      RECT 1052.3500 702.7150 1057.5000 705.7150 ;
      RECT 1044.2000 702.7150 1049.3500 705.7150 ;
      RECT 1036.0500 702.7150 1041.2000 705.7150 ;
      RECT 1027.9000 702.7150 1033.0500 705.7150 ;
      RECT 1019.7500 702.7150 1024.9000 705.7150 ;
      RECT 1011.6000 702.7150 1016.7500 705.7150 ;
      RECT 1003.4500 702.7150 1008.6000 705.7150 ;
      RECT 995.3000 702.7150 1000.4500 705.7150 ;
      RECT 987.1500 702.7150 992.3000 705.7150 ;
      RECT 979.0000 702.7150 984.1500 705.7150 ;
      RECT 970.8500 702.7150 976.0000 705.7150 ;
      RECT 962.7000 702.7150 967.8500 705.7150 ;
      RECT 954.5500 702.7150 959.7000 705.7150 ;
      RECT 946.4000 702.7150 951.5500 705.7150 ;
      RECT 938.2500 702.7150 943.4000 705.7150 ;
      RECT 930.1000 702.7150 935.2500 705.7150 ;
      RECT 921.9500 702.7150 927.1000 705.7150 ;
      RECT 913.8000 702.7150 918.9500 705.7150 ;
      RECT 905.6500 702.7150 910.8000 705.7150 ;
      RECT 897.5000 702.7150 902.6500 705.7150 ;
      RECT 889.3500 702.7150 894.5000 705.7150 ;
      RECT 881.2000 702.7150 886.3500 705.7150 ;
      RECT 873.0500 702.7150 878.2000 705.7150 ;
      RECT 864.9000 702.7150 870.0500 705.7150 ;
      RECT 856.7500 702.7150 861.9000 705.7150 ;
      RECT 848.6000 702.7150 853.7500 705.7150 ;
      RECT 840.4500 702.7150 845.6000 705.7150 ;
      RECT 832.3000 702.7150 837.4500 705.7150 ;
      RECT 824.1500 702.7150 829.3000 705.7150 ;
      RECT 816.0000 702.7150 821.1500 705.7150 ;
      RECT 807.8500 702.7150 813.0000 705.7150 ;
      RECT 799.7000 702.7150 804.8500 705.7150 ;
      RECT 791.5500 702.7150 796.7000 705.7150 ;
      RECT 783.4000 702.7150 788.5500 705.7150 ;
      RECT 775.2500 702.7150 780.4000 705.7150 ;
      RECT 767.1000 702.7150 772.2500 705.7150 ;
      RECT 758.9500 702.7150 764.1000 705.7150 ;
      RECT 750.8000 702.7150 755.9500 705.7150 ;
      RECT 742.6500 702.7150 747.8000 705.7150 ;
      RECT 734.5000 702.7150 739.6500 705.7150 ;
      RECT 726.3500 702.7150 731.5000 705.7150 ;
      RECT 718.2000 702.7150 723.3500 705.7150 ;
      RECT 710.0500 702.7150 715.2000 705.7150 ;
      RECT 701.9000 702.7150 707.0500 705.7150 ;
      RECT 693.7500 702.7150 698.9000 705.7150 ;
      RECT 685.6000 702.7150 690.7500 705.7150 ;
      RECT 677.4500 702.7150 682.6000 705.7150 ;
      RECT 669.3000 702.7150 674.4500 705.7150 ;
      RECT 661.1500 702.7150 666.3000 705.7150 ;
      RECT 653.0000 702.7150 658.1500 705.7150 ;
      RECT 644.8500 702.7150 650.0000 705.7150 ;
      RECT 636.7000 702.7150 641.8500 705.7150 ;
      RECT 628.5500 702.7150 633.7000 705.7150 ;
      RECT 620.4000 702.7150 625.5500 705.7150 ;
      RECT 612.2500 702.7150 617.4000 705.7150 ;
      RECT 604.1000 702.7150 609.2500 705.7150 ;
      RECT 595.9500 702.7150 601.1000 705.7150 ;
      RECT 587.8000 702.7150 592.9500 705.7150 ;
      RECT 579.6500 702.7150 584.8000 705.7150 ;
      RECT 571.5000 702.7150 576.6500 705.7150 ;
      RECT 563.3500 702.7150 568.5000 705.7150 ;
      RECT 555.2000 702.7150 560.3500 705.7150 ;
      RECT 547.0500 702.7150 552.2000 705.7150 ;
      RECT 538.9000 702.7150 544.0500 705.7150 ;
      RECT 530.7500 702.7150 535.9000 705.7150 ;
      RECT 522.6000 702.7150 527.7500 705.7150 ;
      RECT 514.4500 702.7150 519.6000 705.7150 ;
      RECT 506.3000 702.7150 511.4500 705.7150 ;
      RECT 498.1500 702.7150 503.3000 705.7150 ;
      RECT 490.0000 702.7150 495.1500 705.7150 ;
      RECT 481.8500 702.7150 487.0000 705.7150 ;
      RECT 473.7000 702.7150 478.8500 705.7150 ;
      RECT 465.5500 702.7150 470.7000 705.7150 ;
      RECT 457.4000 702.7150 462.5500 705.7150 ;
      RECT 449.2500 702.7150 454.4000 705.7150 ;
      RECT 441.1000 702.7150 446.2500 705.7150 ;
      RECT 432.9500 702.7150 438.1000 705.7150 ;
      RECT 424.8000 702.7150 429.9500 705.7150 ;
      RECT 416.6500 702.7150 421.8000 705.7150 ;
      RECT 396.5000 702.7150 413.6500 705.7150 ;
      RECT 8.5000 702.7150 393.5000 705.7150 ;
      RECT 0.0000 702.7150 5.5000 705.7150 ;
      RECT 0.0000 701.3000 1120.0000 702.7150 ;
      RECT 1116.6000 700.7150 1120.0000 701.3000 ;
      RECT 0.0000 698.6200 1113.6000 701.3000 ;
      RECT 1118.5000 697.7150 1120.0000 700.7150 ;
      RECT 1114.5000 695.6200 1120.0000 697.7150 ;
      RECT 1076.5000 695.6200 1111.5000 698.6200 ;
      RECT 1060.5000 695.6200 1073.5000 698.6200 ;
      RECT 1052.3500 695.6200 1057.5000 698.6200 ;
      RECT 1044.2000 695.6200 1049.3500 698.6200 ;
      RECT 1036.0500 695.6200 1041.2000 698.6200 ;
      RECT 1027.9000 695.6200 1033.0500 698.6200 ;
      RECT 1019.7500 695.6200 1024.9000 698.6200 ;
      RECT 1011.6000 695.6200 1016.7500 698.6200 ;
      RECT 1003.4500 695.6200 1008.6000 698.6200 ;
      RECT 995.3000 695.6200 1000.4500 698.6200 ;
      RECT 987.1500 695.6200 992.3000 698.6200 ;
      RECT 979.0000 695.6200 984.1500 698.6200 ;
      RECT 970.8500 695.6200 976.0000 698.6200 ;
      RECT 962.7000 695.6200 967.8500 698.6200 ;
      RECT 954.5500 695.6200 959.7000 698.6200 ;
      RECT 946.4000 695.6200 951.5500 698.6200 ;
      RECT 938.2500 695.6200 943.4000 698.6200 ;
      RECT 930.1000 695.6200 935.2500 698.6200 ;
      RECT 921.9500 695.6200 927.1000 698.6200 ;
      RECT 913.8000 695.6200 918.9500 698.6200 ;
      RECT 905.6500 695.6200 910.8000 698.6200 ;
      RECT 897.5000 695.6200 902.6500 698.6200 ;
      RECT 889.3500 695.6200 894.5000 698.6200 ;
      RECT 881.2000 695.6200 886.3500 698.6200 ;
      RECT 873.0500 695.6200 878.2000 698.6200 ;
      RECT 864.9000 695.6200 870.0500 698.6200 ;
      RECT 856.7500 695.6200 861.9000 698.6200 ;
      RECT 848.6000 695.6200 853.7500 698.6200 ;
      RECT 840.4500 695.6200 845.6000 698.6200 ;
      RECT 832.3000 695.6200 837.4500 698.6200 ;
      RECT 824.1500 695.6200 829.3000 698.6200 ;
      RECT 816.0000 695.6200 821.1500 698.6200 ;
      RECT 807.8500 695.6200 813.0000 698.6200 ;
      RECT 799.7000 695.6200 804.8500 698.6200 ;
      RECT 791.5500 695.6200 796.7000 698.6200 ;
      RECT 783.4000 695.6200 788.5500 698.6200 ;
      RECT 775.2500 695.6200 780.4000 698.6200 ;
      RECT 767.1000 695.6200 772.2500 698.6200 ;
      RECT 758.9500 695.6200 764.1000 698.6200 ;
      RECT 750.8000 695.6200 755.9500 698.6200 ;
      RECT 742.6500 695.6200 747.8000 698.6200 ;
      RECT 734.5000 695.6200 739.6500 698.6200 ;
      RECT 726.3500 695.6200 731.5000 698.6200 ;
      RECT 718.2000 695.6200 723.3500 698.6200 ;
      RECT 710.0500 695.6200 715.2000 698.6200 ;
      RECT 701.9000 695.6200 707.0500 698.6200 ;
      RECT 693.7500 695.6200 698.9000 698.6200 ;
      RECT 685.6000 695.6200 690.7500 698.6200 ;
      RECT 677.4500 695.6200 682.6000 698.6200 ;
      RECT 669.3000 695.6200 674.4500 698.6200 ;
      RECT 661.1500 695.6200 666.3000 698.6200 ;
      RECT 653.0000 695.6200 658.1500 698.6200 ;
      RECT 644.8500 695.6200 650.0000 698.6200 ;
      RECT 636.7000 695.6200 641.8500 698.6200 ;
      RECT 628.5500 695.6200 633.7000 698.6200 ;
      RECT 620.4000 695.6200 625.5500 698.6200 ;
      RECT 612.2500 695.6200 617.4000 698.6200 ;
      RECT 604.1000 695.6200 609.2500 698.6200 ;
      RECT 595.9500 695.6200 601.1000 698.6200 ;
      RECT 587.8000 695.6200 592.9500 698.6200 ;
      RECT 579.6500 695.6200 584.8000 698.6200 ;
      RECT 571.5000 695.6200 576.6500 698.6200 ;
      RECT 563.3500 695.6200 568.5000 698.6200 ;
      RECT 555.2000 695.6200 560.3500 698.6200 ;
      RECT 547.0500 695.6200 552.2000 698.6200 ;
      RECT 538.9000 695.6200 544.0500 698.6200 ;
      RECT 530.7500 695.6200 535.9000 698.6200 ;
      RECT 522.6000 695.6200 527.7500 698.6200 ;
      RECT 514.4500 695.6200 519.6000 698.6200 ;
      RECT 506.3000 695.6200 511.4500 698.6200 ;
      RECT 498.1500 695.6200 503.3000 698.6200 ;
      RECT 490.0000 695.6200 495.1500 698.6200 ;
      RECT 481.8500 695.6200 487.0000 698.6200 ;
      RECT 473.7000 695.6200 478.8500 698.6200 ;
      RECT 465.5500 695.6200 470.7000 698.6200 ;
      RECT 457.4000 695.6200 462.5500 698.6200 ;
      RECT 449.2500 695.6200 454.4000 698.6200 ;
      RECT 441.1000 695.6200 446.2500 698.6200 ;
      RECT 432.9500 695.6200 438.1000 698.6200 ;
      RECT 424.8000 695.6200 429.9500 698.6200 ;
      RECT 416.6500 695.6200 421.8000 698.6200 ;
      RECT 396.5000 695.6200 413.6500 698.6200 ;
      RECT 8.5000 695.6200 393.5000 698.6200 ;
      RECT 0.0000 695.6200 5.5000 698.6200 ;
      RECT 0.0000 694.1000 1120.0000 695.6200 ;
      RECT 1116.6000 693.6200 1120.0000 694.1000 ;
      RECT 0.0000 693.5000 1113.6000 694.1000 ;
      RECT 330.4650 691.5250 1113.6000 693.5000 ;
      RECT 0.0000 691.5250 327.4650 693.5000 ;
      RECT 330.4650 691.0250 343.5000 691.5250 ;
      RECT 46.5000 691.0250 327.4650 691.5250 ;
      RECT 1118.5000 690.6200 1120.0000 693.6200 ;
      RECT 1114.5000 688.5250 1120.0000 690.6200 ;
      RECT 1076.5000 688.5250 1111.5000 691.5250 ;
      RECT 1060.5000 688.5250 1073.5000 691.5250 ;
      RECT 1052.3500 688.5250 1057.5000 691.5250 ;
      RECT 1044.2000 688.5250 1049.3500 691.5250 ;
      RECT 1036.0500 688.5250 1041.2000 691.5250 ;
      RECT 1027.9000 688.5250 1033.0500 691.5250 ;
      RECT 1019.7500 688.5250 1024.9000 691.5250 ;
      RECT 1011.6000 688.5250 1016.7500 691.5250 ;
      RECT 1003.4500 688.5250 1008.6000 691.5250 ;
      RECT 995.3000 688.5250 1000.4500 691.5250 ;
      RECT 987.1500 688.5250 992.3000 691.5250 ;
      RECT 979.0000 688.5250 984.1500 691.5250 ;
      RECT 970.8500 688.5250 976.0000 691.5250 ;
      RECT 962.7000 688.5250 967.8500 691.5250 ;
      RECT 954.5500 688.5250 959.7000 691.5250 ;
      RECT 946.4000 688.5250 951.5500 691.5250 ;
      RECT 938.2500 688.5250 943.4000 691.5250 ;
      RECT 930.1000 688.5250 935.2500 691.5250 ;
      RECT 921.9500 688.5250 927.1000 691.5250 ;
      RECT 913.8000 688.5250 918.9500 691.5250 ;
      RECT 905.6500 688.5250 910.8000 691.5250 ;
      RECT 897.5000 688.5250 902.6500 691.5250 ;
      RECT 889.3500 688.5250 894.5000 691.5250 ;
      RECT 881.2000 688.5250 886.3500 691.5250 ;
      RECT 873.0500 688.5250 878.2000 691.5250 ;
      RECT 864.9000 688.5250 870.0500 691.5250 ;
      RECT 856.7500 688.5250 861.9000 691.5250 ;
      RECT 848.6000 688.5250 853.7500 691.5250 ;
      RECT 840.4500 688.5250 845.6000 691.5250 ;
      RECT 832.3000 688.5250 837.4500 691.5250 ;
      RECT 824.1500 688.5250 829.3000 691.5250 ;
      RECT 816.0000 688.5250 821.1500 691.5250 ;
      RECT 807.8500 688.5250 813.0000 691.5250 ;
      RECT 799.7000 688.5250 804.8500 691.5250 ;
      RECT 791.5500 688.5250 796.7000 691.5250 ;
      RECT 783.4000 688.5250 788.5500 691.5250 ;
      RECT 775.2500 688.5250 780.4000 691.5250 ;
      RECT 767.1000 688.5250 772.2500 691.5250 ;
      RECT 758.9500 688.5250 764.1000 691.5250 ;
      RECT 750.8000 688.5250 755.9500 691.5250 ;
      RECT 742.6500 688.5250 747.8000 691.5250 ;
      RECT 734.5000 688.5250 739.6500 691.5250 ;
      RECT 726.3500 688.5250 731.5000 691.5250 ;
      RECT 718.2000 688.5250 723.3500 691.5250 ;
      RECT 710.0500 688.5250 715.2000 691.5250 ;
      RECT 701.9000 688.5250 707.0500 691.5250 ;
      RECT 693.7500 688.5250 698.9000 691.5250 ;
      RECT 685.6000 688.5250 690.7500 691.5250 ;
      RECT 677.4500 688.5250 682.6000 691.5250 ;
      RECT 669.3000 688.5250 674.4500 691.5250 ;
      RECT 661.1500 688.5250 666.3000 691.5250 ;
      RECT 653.0000 688.5250 658.1500 691.5250 ;
      RECT 644.8500 688.5250 650.0000 691.5250 ;
      RECT 636.7000 688.5250 641.8500 691.5250 ;
      RECT 628.5500 688.5250 633.7000 691.5250 ;
      RECT 620.4000 688.5250 625.5500 691.5250 ;
      RECT 612.2500 688.5250 617.4000 691.5250 ;
      RECT 604.1000 688.5250 609.2500 691.5250 ;
      RECT 595.9500 688.5250 601.1000 691.5250 ;
      RECT 587.8000 688.5250 592.9500 691.5250 ;
      RECT 579.6500 688.5250 584.8000 691.5250 ;
      RECT 571.5000 688.5250 576.6500 691.5250 ;
      RECT 563.3500 688.5250 568.5000 691.5250 ;
      RECT 555.2000 688.5250 560.3500 691.5250 ;
      RECT 547.0500 688.5250 552.2000 691.5250 ;
      RECT 538.9000 688.5250 544.0500 691.5250 ;
      RECT 530.7500 688.5250 535.9000 691.5250 ;
      RECT 522.6000 688.5250 527.7500 691.5250 ;
      RECT 514.4500 688.5250 519.6000 691.5250 ;
      RECT 506.3000 688.5250 511.4500 691.5250 ;
      RECT 498.1500 688.5250 503.3000 691.5250 ;
      RECT 490.0000 688.5250 495.1500 691.5250 ;
      RECT 481.8500 688.5250 487.0000 691.5250 ;
      RECT 473.7000 688.5250 478.8500 691.5250 ;
      RECT 465.5500 688.5250 470.7000 691.5250 ;
      RECT 457.4000 688.5250 462.5500 691.5250 ;
      RECT 449.2500 688.5250 454.4000 691.5250 ;
      RECT 441.1000 688.5250 446.2500 691.5250 ;
      RECT 432.9500 688.5250 438.1000 691.5250 ;
      RECT 424.8000 688.5250 429.9500 691.5250 ;
      RECT 416.6500 688.5250 421.8000 691.5250 ;
      RECT 396.5000 688.5250 413.6500 691.5250 ;
      RECT 346.5000 688.5250 393.5000 691.5250 ;
      RECT 46.5000 688.5250 343.5000 691.0250 ;
      RECT 8.5000 688.5250 43.5000 691.5250 ;
      RECT 0.0000 688.5250 5.5000 691.5250 ;
      RECT 0.0000 687.1000 1120.0000 688.5250 ;
      RECT 1116.6000 686.5250 1120.0000 687.1000 ;
      RECT 0.0000 684.4300 1113.6000 687.1000 ;
      RECT 1118.5000 683.5250 1120.0000 686.5250 ;
      RECT 1114.5000 681.4300 1120.0000 683.5250 ;
      RECT 1076.5000 681.4300 1111.5000 684.4300 ;
      RECT 1060.5000 681.4300 1073.5000 684.4300 ;
      RECT 1052.3500 681.4300 1057.5000 684.4300 ;
      RECT 1044.2000 681.4300 1049.3500 684.4300 ;
      RECT 1036.0500 681.4300 1041.2000 684.4300 ;
      RECT 1027.9000 681.4300 1033.0500 684.4300 ;
      RECT 1019.7500 681.4300 1024.9000 684.4300 ;
      RECT 1011.6000 681.4300 1016.7500 684.4300 ;
      RECT 1003.4500 681.4300 1008.6000 684.4300 ;
      RECT 995.3000 681.4300 1000.4500 684.4300 ;
      RECT 987.1500 681.4300 992.3000 684.4300 ;
      RECT 979.0000 681.4300 984.1500 684.4300 ;
      RECT 970.8500 681.4300 976.0000 684.4300 ;
      RECT 962.7000 681.4300 967.8500 684.4300 ;
      RECT 954.5500 681.4300 959.7000 684.4300 ;
      RECT 946.4000 681.4300 951.5500 684.4300 ;
      RECT 938.2500 681.4300 943.4000 684.4300 ;
      RECT 930.1000 681.4300 935.2500 684.4300 ;
      RECT 921.9500 681.4300 927.1000 684.4300 ;
      RECT 913.8000 681.4300 918.9500 684.4300 ;
      RECT 905.6500 681.4300 910.8000 684.4300 ;
      RECT 897.5000 681.4300 902.6500 684.4300 ;
      RECT 889.3500 681.4300 894.5000 684.4300 ;
      RECT 881.2000 681.4300 886.3500 684.4300 ;
      RECT 873.0500 681.4300 878.2000 684.4300 ;
      RECT 864.9000 681.4300 870.0500 684.4300 ;
      RECT 856.7500 681.4300 861.9000 684.4300 ;
      RECT 848.6000 681.4300 853.7500 684.4300 ;
      RECT 840.4500 681.4300 845.6000 684.4300 ;
      RECT 832.3000 681.4300 837.4500 684.4300 ;
      RECT 824.1500 681.4300 829.3000 684.4300 ;
      RECT 816.0000 681.4300 821.1500 684.4300 ;
      RECT 807.8500 681.4300 813.0000 684.4300 ;
      RECT 799.7000 681.4300 804.8500 684.4300 ;
      RECT 791.5500 681.4300 796.7000 684.4300 ;
      RECT 783.4000 681.4300 788.5500 684.4300 ;
      RECT 775.2500 681.4300 780.4000 684.4300 ;
      RECT 767.1000 681.4300 772.2500 684.4300 ;
      RECT 758.9500 681.4300 764.1000 684.4300 ;
      RECT 750.8000 681.4300 755.9500 684.4300 ;
      RECT 742.6500 681.4300 747.8000 684.4300 ;
      RECT 734.5000 681.4300 739.6500 684.4300 ;
      RECT 726.3500 681.4300 731.5000 684.4300 ;
      RECT 718.2000 681.4300 723.3500 684.4300 ;
      RECT 710.0500 681.4300 715.2000 684.4300 ;
      RECT 701.9000 681.4300 707.0500 684.4300 ;
      RECT 693.7500 681.4300 698.9000 684.4300 ;
      RECT 685.6000 681.4300 690.7500 684.4300 ;
      RECT 677.4500 681.4300 682.6000 684.4300 ;
      RECT 669.3000 681.4300 674.4500 684.4300 ;
      RECT 661.1500 681.4300 666.3000 684.4300 ;
      RECT 653.0000 681.4300 658.1500 684.4300 ;
      RECT 644.8500 681.4300 650.0000 684.4300 ;
      RECT 636.7000 681.4300 641.8500 684.4300 ;
      RECT 628.5500 681.4300 633.7000 684.4300 ;
      RECT 620.4000 681.4300 625.5500 684.4300 ;
      RECT 612.2500 681.4300 617.4000 684.4300 ;
      RECT 604.1000 681.4300 609.2500 684.4300 ;
      RECT 595.9500 681.4300 601.1000 684.4300 ;
      RECT 587.8000 681.4300 592.9500 684.4300 ;
      RECT 579.6500 681.4300 584.8000 684.4300 ;
      RECT 571.5000 681.4300 576.6500 684.4300 ;
      RECT 563.3500 681.4300 568.5000 684.4300 ;
      RECT 555.2000 681.4300 560.3500 684.4300 ;
      RECT 547.0500 681.4300 552.2000 684.4300 ;
      RECT 538.9000 681.4300 544.0500 684.4300 ;
      RECT 530.7500 681.4300 535.9000 684.4300 ;
      RECT 522.6000 681.4300 527.7500 684.4300 ;
      RECT 514.4500 681.4300 519.6000 684.4300 ;
      RECT 506.3000 681.4300 511.4500 684.4300 ;
      RECT 498.1500 681.4300 503.3000 684.4300 ;
      RECT 490.0000 681.4300 495.1500 684.4300 ;
      RECT 481.8500 681.4300 487.0000 684.4300 ;
      RECT 473.7000 681.4300 478.8500 684.4300 ;
      RECT 465.5500 681.4300 470.7000 684.4300 ;
      RECT 457.4000 681.4300 462.5500 684.4300 ;
      RECT 449.2500 681.4300 454.4000 684.4300 ;
      RECT 441.1000 681.4300 446.2500 684.4300 ;
      RECT 432.9500 681.4300 438.1000 684.4300 ;
      RECT 424.8000 681.4300 429.9500 684.4300 ;
      RECT 416.6500 681.4300 421.8000 684.4300 ;
      RECT 396.5000 681.4300 413.6500 684.4300 ;
      RECT 346.5000 681.4300 393.5000 684.4300 ;
      RECT 46.5000 681.4300 343.5000 684.4300 ;
      RECT 8.5000 681.4300 43.5000 684.4300 ;
      RECT 0.0000 681.4300 5.5000 684.4300 ;
      RECT 0.0000 680.5000 1120.0000 681.4300 ;
      RECT 62.5000 679.9000 1120.0000 680.5000 ;
      RECT 62.5000 679.8350 1113.6000 679.9000 ;
      RECT 1116.6000 679.4300 1120.0000 679.9000 ;
      RECT 330.4650 677.6650 1113.6000 679.8350 ;
      RECT 62.5000 677.6650 327.4650 679.8350 ;
      RECT 62.5000 677.5000 1113.6000 677.6650 ;
      RECT 0.0000 677.5000 59.5000 680.5000 ;
      RECT 0.0000 677.3350 1113.6000 677.5000 ;
      RECT 1118.5000 676.4300 1120.0000 679.4300 ;
      RECT 1114.5000 674.3350 1120.0000 676.4300 ;
      RECT 1076.5000 674.3350 1111.5000 677.3350 ;
      RECT 1060.5000 674.3350 1073.5000 677.3350 ;
      RECT 1052.3500 674.3350 1057.5000 677.3350 ;
      RECT 1044.2000 674.3350 1049.3500 677.3350 ;
      RECT 1036.0500 674.3350 1041.2000 677.3350 ;
      RECT 1027.9000 674.3350 1033.0500 677.3350 ;
      RECT 1019.7500 674.3350 1024.9000 677.3350 ;
      RECT 1011.6000 674.3350 1016.7500 677.3350 ;
      RECT 1003.4500 674.3350 1008.6000 677.3350 ;
      RECT 995.3000 674.3350 1000.4500 677.3350 ;
      RECT 987.1500 674.3350 992.3000 677.3350 ;
      RECT 979.0000 674.3350 984.1500 677.3350 ;
      RECT 970.8500 674.3350 976.0000 677.3350 ;
      RECT 962.7000 674.3350 967.8500 677.3350 ;
      RECT 954.5500 674.3350 959.7000 677.3350 ;
      RECT 946.4000 674.3350 951.5500 677.3350 ;
      RECT 938.2500 674.3350 943.4000 677.3350 ;
      RECT 930.1000 674.3350 935.2500 677.3350 ;
      RECT 921.9500 674.3350 927.1000 677.3350 ;
      RECT 913.8000 674.3350 918.9500 677.3350 ;
      RECT 905.6500 674.3350 910.8000 677.3350 ;
      RECT 897.5000 674.3350 902.6500 677.3350 ;
      RECT 889.3500 674.3350 894.5000 677.3350 ;
      RECT 881.2000 674.3350 886.3500 677.3350 ;
      RECT 873.0500 674.3350 878.2000 677.3350 ;
      RECT 864.9000 674.3350 870.0500 677.3350 ;
      RECT 856.7500 674.3350 861.9000 677.3350 ;
      RECT 848.6000 674.3350 853.7500 677.3350 ;
      RECT 840.4500 674.3350 845.6000 677.3350 ;
      RECT 832.3000 674.3350 837.4500 677.3350 ;
      RECT 824.1500 674.3350 829.3000 677.3350 ;
      RECT 816.0000 674.3350 821.1500 677.3350 ;
      RECT 807.8500 674.3350 813.0000 677.3350 ;
      RECT 799.7000 674.3350 804.8500 677.3350 ;
      RECT 791.5500 674.3350 796.7000 677.3350 ;
      RECT 783.4000 674.3350 788.5500 677.3350 ;
      RECT 775.2500 674.3350 780.4000 677.3350 ;
      RECT 767.1000 674.3350 772.2500 677.3350 ;
      RECT 758.9500 674.3350 764.1000 677.3350 ;
      RECT 750.8000 674.3350 755.9500 677.3350 ;
      RECT 742.6500 674.3350 747.8000 677.3350 ;
      RECT 734.5000 674.3350 739.6500 677.3350 ;
      RECT 726.3500 674.3350 731.5000 677.3350 ;
      RECT 718.2000 674.3350 723.3500 677.3350 ;
      RECT 710.0500 674.3350 715.2000 677.3350 ;
      RECT 701.9000 674.3350 707.0500 677.3350 ;
      RECT 693.7500 674.3350 698.9000 677.3350 ;
      RECT 685.6000 674.3350 690.7500 677.3350 ;
      RECT 677.4500 674.3350 682.6000 677.3350 ;
      RECT 669.3000 674.3350 674.4500 677.3350 ;
      RECT 661.1500 674.3350 666.3000 677.3350 ;
      RECT 653.0000 674.3350 658.1500 677.3350 ;
      RECT 644.8500 674.3350 650.0000 677.3350 ;
      RECT 636.7000 674.3350 641.8500 677.3350 ;
      RECT 628.5500 674.3350 633.7000 677.3350 ;
      RECT 620.4000 674.3350 625.5500 677.3350 ;
      RECT 612.2500 674.3350 617.4000 677.3350 ;
      RECT 604.1000 674.3350 609.2500 677.3350 ;
      RECT 595.9500 674.3350 601.1000 677.3350 ;
      RECT 587.8000 674.3350 592.9500 677.3350 ;
      RECT 579.6500 674.3350 584.8000 677.3350 ;
      RECT 571.5000 674.3350 576.6500 677.3350 ;
      RECT 563.3500 674.3350 568.5000 677.3350 ;
      RECT 555.2000 674.3350 560.3500 677.3350 ;
      RECT 547.0500 674.3350 552.2000 677.3350 ;
      RECT 538.9000 674.3350 544.0500 677.3350 ;
      RECT 530.7500 674.3350 535.9000 677.3350 ;
      RECT 522.6000 674.3350 527.7500 677.3350 ;
      RECT 514.4500 674.3350 519.6000 677.3350 ;
      RECT 506.3000 674.3350 511.4500 677.3350 ;
      RECT 498.1500 674.3350 503.3000 677.3350 ;
      RECT 490.0000 674.3350 495.1500 677.3350 ;
      RECT 481.8500 674.3350 487.0000 677.3350 ;
      RECT 473.7000 674.3350 478.8500 677.3350 ;
      RECT 465.5500 674.3350 470.7000 677.3350 ;
      RECT 457.4000 674.3350 462.5500 677.3350 ;
      RECT 449.2500 674.3350 454.4000 677.3350 ;
      RECT 441.1000 674.3350 446.2500 677.3350 ;
      RECT 432.9500 674.3350 438.1000 677.3350 ;
      RECT 424.8000 674.3350 429.9500 677.3350 ;
      RECT 416.6500 674.3350 421.8000 677.3350 ;
      RECT 396.5000 674.3350 413.6500 677.3350 ;
      RECT 346.5000 674.3350 393.5000 677.3350 ;
      RECT 326.4650 674.3350 343.5000 677.3350 ;
      RECT 317.9500 674.3350 323.4650 677.3350 ;
      RECT 309.4350 674.3350 314.9500 677.3350 ;
      RECT 300.9200 674.3350 306.4350 677.3350 ;
      RECT 292.4050 674.3350 297.9200 677.3350 ;
      RECT 283.8900 674.3350 289.4050 677.3350 ;
      RECT 275.3750 674.3350 280.8900 677.3350 ;
      RECT 266.8600 674.3350 272.3750 677.3350 ;
      RECT 258.3450 674.3350 263.8600 677.3350 ;
      RECT 249.8300 674.3350 255.3450 677.3350 ;
      RECT 241.3150 674.3350 246.8300 677.3350 ;
      RECT 232.8000 674.3350 238.3150 677.3350 ;
      RECT 224.2850 674.3350 229.8000 677.3350 ;
      RECT 215.7700 674.3350 221.2850 677.3350 ;
      RECT 207.2550 674.3350 212.7700 677.3350 ;
      RECT 198.7400 674.3350 204.2550 677.3350 ;
      RECT 190.2250 674.3350 195.7400 677.3350 ;
      RECT 181.7100 674.3350 187.2250 677.3350 ;
      RECT 173.1950 674.3350 178.7100 677.3350 ;
      RECT 164.6800 674.3350 170.1950 677.3350 ;
      RECT 156.1650 674.3350 161.6800 677.3350 ;
      RECT 147.6500 674.3350 153.1650 677.3350 ;
      RECT 139.1350 674.3350 144.6500 677.3350 ;
      RECT 130.6200 674.3350 136.1350 677.3350 ;
      RECT 122.1050 674.3350 127.6200 677.3350 ;
      RECT 113.5900 674.3350 119.1050 677.3350 ;
      RECT 105.0750 674.3350 110.5900 677.3350 ;
      RECT 96.5600 674.3350 102.0750 677.3350 ;
      RECT 88.0450 674.3350 93.5600 677.3350 ;
      RECT 79.5300 674.3350 85.0450 677.3350 ;
      RECT 71.0150 674.3350 76.5300 677.3350 ;
      RECT 62.5000 674.3350 68.0150 677.3350 ;
      RECT 46.5000 674.3350 59.5000 677.3350 ;
      RECT 8.5000 674.3350 43.5000 677.3350 ;
      RECT 0.0000 674.3350 5.5000 677.3350 ;
      RECT 0.0000 672.9000 1120.0000 674.3350 ;
      RECT 1116.6000 672.3350 1120.0000 672.9000 ;
      RECT 0.0000 670.2400 1113.6000 672.9000 ;
      RECT 1118.5000 669.3350 1120.0000 672.3350 ;
      RECT 1114.5000 667.2400 1120.0000 669.3350 ;
      RECT 1076.5000 667.2400 1111.5000 670.2400 ;
      RECT 1060.5000 667.2400 1073.5000 670.2400 ;
      RECT 1052.3500 667.2400 1057.5000 670.2400 ;
      RECT 1044.2000 667.2400 1049.3500 670.2400 ;
      RECT 1036.0500 667.2400 1041.2000 670.2400 ;
      RECT 1027.9000 667.2400 1033.0500 670.2400 ;
      RECT 1019.7500 667.2400 1024.9000 670.2400 ;
      RECT 1011.6000 667.2400 1016.7500 670.2400 ;
      RECT 1003.4500 667.2400 1008.6000 670.2400 ;
      RECT 995.3000 667.2400 1000.4500 670.2400 ;
      RECT 987.1500 667.2400 992.3000 670.2400 ;
      RECT 979.0000 667.2400 984.1500 670.2400 ;
      RECT 970.8500 667.2400 976.0000 670.2400 ;
      RECT 962.7000 667.2400 967.8500 670.2400 ;
      RECT 954.5500 667.2400 959.7000 670.2400 ;
      RECT 946.4000 667.2400 951.5500 670.2400 ;
      RECT 938.2500 667.2400 943.4000 670.2400 ;
      RECT 930.1000 667.2400 935.2500 670.2400 ;
      RECT 921.9500 667.2400 927.1000 670.2400 ;
      RECT 913.8000 667.2400 918.9500 670.2400 ;
      RECT 905.6500 667.2400 910.8000 670.2400 ;
      RECT 897.5000 667.2400 902.6500 670.2400 ;
      RECT 889.3500 667.2400 894.5000 670.2400 ;
      RECT 881.2000 667.2400 886.3500 670.2400 ;
      RECT 873.0500 667.2400 878.2000 670.2400 ;
      RECT 864.9000 667.2400 870.0500 670.2400 ;
      RECT 856.7500 667.2400 861.9000 670.2400 ;
      RECT 848.6000 667.2400 853.7500 670.2400 ;
      RECT 840.4500 667.2400 845.6000 670.2400 ;
      RECT 832.3000 667.2400 837.4500 670.2400 ;
      RECT 824.1500 667.2400 829.3000 670.2400 ;
      RECT 816.0000 667.2400 821.1500 670.2400 ;
      RECT 807.8500 667.2400 813.0000 670.2400 ;
      RECT 799.7000 667.2400 804.8500 670.2400 ;
      RECT 791.5500 667.2400 796.7000 670.2400 ;
      RECT 783.4000 667.2400 788.5500 670.2400 ;
      RECT 775.2500 667.2400 780.4000 670.2400 ;
      RECT 767.1000 667.2400 772.2500 670.2400 ;
      RECT 758.9500 667.2400 764.1000 670.2400 ;
      RECT 750.8000 667.2400 755.9500 670.2400 ;
      RECT 742.6500 667.2400 747.8000 670.2400 ;
      RECT 734.5000 667.2400 739.6500 670.2400 ;
      RECT 726.3500 667.2400 731.5000 670.2400 ;
      RECT 718.2000 667.2400 723.3500 670.2400 ;
      RECT 710.0500 667.2400 715.2000 670.2400 ;
      RECT 701.9000 667.2400 707.0500 670.2400 ;
      RECT 693.7500 667.2400 698.9000 670.2400 ;
      RECT 685.6000 667.2400 690.7500 670.2400 ;
      RECT 677.4500 667.2400 682.6000 670.2400 ;
      RECT 669.3000 667.2400 674.4500 670.2400 ;
      RECT 661.1500 667.2400 666.3000 670.2400 ;
      RECT 653.0000 667.2400 658.1500 670.2400 ;
      RECT 644.8500 667.2400 650.0000 670.2400 ;
      RECT 636.7000 667.2400 641.8500 670.2400 ;
      RECT 628.5500 667.2400 633.7000 670.2400 ;
      RECT 620.4000 667.2400 625.5500 670.2400 ;
      RECT 612.2500 667.2400 617.4000 670.2400 ;
      RECT 604.1000 667.2400 609.2500 670.2400 ;
      RECT 595.9500 667.2400 601.1000 670.2400 ;
      RECT 587.8000 667.2400 592.9500 670.2400 ;
      RECT 579.6500 667.2400 584.8000 670.2400 ;
      RECT 571.5000 667.2400 576.6500 670.2400 ;
      RECT 563.3500 667.2400 568.5000 670.2400 ;
      RECT 555.2000 667.2400 560.3500 670.2400 ;
      RECT 547.0500 667.2400 552.2000 670.2400 ;
      RECT 538.9000 667.2400 544.0500 670.2400 ;
      RECT 530.7500 667.2400 535.9000 670.2400 ;
      RECT 522.6000 667.2400 527.7500 670.2400 ;
      RECT 514.4500 667.2400 519.6000 670.2400 ;
      RECT 506.3000 667.2400 511.4500 670.2400 ;
      RECT 498.1500 667.2400 503.3000 670.2400 ;
      RECT 490.0000 667.2400 495.1500 670.2400 ;
      RECT 481.8500 667.2400 487.0000 670.2400 ;
      RECT 473.7000 667.2400 478.8500 670.2400 ;
      RECT 465.5500 667.2400 470.7000 670.2400 ;
      RECT 457.4000 667.2400 462.5500 670.2400 ;
      RECT 449.2500 667.2400 454.4000 670.2400 ;
      RECT 441.1000 667.2400 446.2500 670.2400 ;
      RECT 432.9500 667.2400 438.1000 670.2400 ;
      RECT 424.8000 667.2400 429.9500 670.2400 ;
      RECT 416.6500 667.2400 421.8000 670.2400 ;
      RECT 396.5000 667.2400 413.6500 670.2400 ;
      RECT 346.5000 667.2400 393.5000 670.2400 ;
      RECT 326.4650 667.2400 343.5000 670.2400 ;
      RECT 317.9500 667.2400 323.4650 670.2400 ;
      RECT 309.4350 667.2400 314.9500 670.2400 ;
      RECT 300.9200 667.2400 306.4350 670.2400 ;
      RECT 292.4050 667.2400 297.9200 670.2400 ;
      RECT 283.8900 667.2400 289.4050 670.2400 ;
      RECT 275.3750 667.2400 280.8900 670.2400 ;
      RECT 266.8600 667.2400 272.3750 670.2400 ;
      RECT 258.3450 667.2400 263.8600 670.2400 ;
      RECT 249.8300 667.2400 255.3450 670.2400 ;
      RECT 241.3150 667.2400 246.8300 670.2400 ;
      RECT 232.8000 667.2400 238.3150 670.2400 ;
      RECT 224.2850 667.2400 229.8000 670.2400 ;
      RECT 215.7700 667.2400 221.2850 670.2400 ;
      RECT 207.2550 667.2400 212.7700 670.2400 ;
      RECT 198.7400 667.2400 204.2550 670.2400 ;
      RECT 190.2250 667.2400 195.7400 670.2400 ;
      RECT 181.7100 667.2400 187.2250 670.2400 ;
      RECT 173.1950 667.2400 178.7100 670.2400 ;
      RECT 164.6800 667.2400 170.1950 670.2400 ;
      RECT 156.1650 667.2400 161.6800 670.2400 ;
      RECT 147.6500 667.2400 153.1650 670.2400 ;
      RECT 139.1350 667.2400 144.6500 670.2400 ;
      RECT 130.6200 667.2400 136.1350 670.2400 ;
      RECT 122.1050 667.2400 127.6200 670.2400 ;
      RECT 113.5900 667.2400 119.1050 670.2400 ;
      RECT 105.0750 667.2400 110.5900 670.2400 ;
      RECT 96.5600 667.2400 102.0750 670.2400 ;
      RECT 88.0450 667.2400 93.5600 670.2400 ;
      RECT 79.5300 667.2400 85.0450 670.2400 ;
      RECT 71.0150 667.2400 76.5300 670.2400 ;
      RECT 62.5000 667.2400 68.0150 670.2400 ;
      RECT 46.5000 667.2400 59.5000 670.2400 ;
      RECT 8.5000 667.2400 43.5000 670.2400 ;
      RECT 0.0000 667.2400 5.5000 670.2400 ;
      RECT 0.0000 665.7000 1120.0000 667.2400 ;
      RECT 1116.6000 665.2400 1120.0000 665.7000 ;
      RECT 0.0000 663.1450 1113.6000 665.7000 ;
      RECT 1118.5000 662.2400 1120.0000 665.2400 ;
      RECT 1114.5000 660.1450 1120.0000 662.2400 ;
      RECT 1076.5000 660.1450 1111.5000 663.1450 ;
      RECT 1060.5000 660.1450 1073.5000 663.1450 ;
      RECT 1052.3500 660.1450 1057.5000 663.1450 ;
      RECT 1044.2000 660.1450 1049.3500 663.1450 ;
      RECT 1036.0500 660.1450 1041.2000 663.1450 ;
      RECT 1027.9000 660.1450 1033.0500 663.1450 ;
      RECT 1019.7500 660.1450 1024.9000 663.1450 ;
      RECT 1011.6000 660.1450 1016.7500 663.1450 ;
      RECT 1003.4500 660.1450 1008.6000 663.1450 ;
      RECT 995.3000 660.1450 1000.4500 663.1450 ;
      RECT 987.1500 660.1450 992.3000 663.1450 ;
      RECT 979.0000 660.1450 984.1500 663.1450 ;
      RECT 970.8500 660.1450 976.0000 663.1450 ;
      RECT 962.7000 660.1450 967.8500 663.1450 ;
      RECT 954.5500 660.1450 959.7000 663.1450 ;
      RECT 946.4000 660.1450 951.5500 663.1450 ;
      RECT 938.2500 660.1450 943.4000 663.1450 ;
      RECT 930.1000 660.1450 935.2500 663.1450 ;
      RECT 921.9500 660.1450 927.1000 663.1450 ;
      RECT 913.8000 660.1450 918.9500 663.1450 ;
      RECT 905.6500 660.1450 910.8000 663.1450 ;
      RECT 897.5000 660.1450 902.6500 663.1450 ;
      RECT 889.3500 660.1450 894.5000 663.1450 ;
      RECT 881.2000 660.1450 886.3500 663.1450 ;
      RECT 873.0500 660.1450 878.2000 663.1450 ;
      RECT 864.9000 660.1450 870.0500 663.1450 ;
      RECT 856.7500 660.1450 861.9000 663.1450 ;
      RECT 848.6000 660.1450 853.7500 663.1450 ;
      RECT 840.4500 660.1450 845.6000 663.1450 ;
      RECT 832.3000 660.1450 837.4500 663.1450 ;
      RECT 824.1500 660.1450 829.3000 663.1450 ;
      RECT 816.0000 660.1450 821.1500 663.1450 ;
      RECT 807.8500 660.1450 813.0000 663.1450 ;
      RECT 799.7000 660.1450 804.8500 663.1450 ;
      RECT 791.5500 660.1450 796.7000 663.1450 ;
      RECT 783.4000 660.1450 788.5500 663.1450 ;
      RECT 775.2500 660.1450 780.4000 663.1450 ;
      RECT 767.1000 660.1450 772.2500 663.1450 ;
      RECT 758.9500 660.1450 764.1000 663.1450 ;
      RECT 750.8000 660.1450 755.9500 663.1450 ;
      RECT 742.6500 660.1450 747.8000 663.1450 ;
      RECT 734.5000 660.1450 739.6500 663.1450 ;
      RECT 726.3500 660.1450 731.5000 663.1450 ;
      RECT 718.2000 660.1450 723.3500 663.1450 ;
      RECT 710.0500 660.1450 715.2000 663.1450 ;
      RECT 701.9000 660.1450 707.0500 663.1450 ;
      RECT 693.7500 660.1450 698.9000 663.1450 ;
      RECT 685.6000 660.1450 690.7500 663.1450 ;
      RECT 677.4500 660.1450 682.6000 663.1450 ;
      RECT 669.3000 660.1450 674.4500 663.1450 ;
      RECT 661.1500 660.1450 666.3000 663.1450 ;
      RECT 653.0000 660.1450 658.1500 663.1450 ;
      RECT 644.8500 660.1450 650.0000 663.1450 ;
      RECT 636.7000 660.1450 641.8500 663.1450 ;
      RECT 628.5500 660.1450 633.7000 663.1450 ;
      RECT 620.4000 660.1450 625.5500 663.1450 ;
      RECT 612.2500 660.1450 617.4000 663.1450 ;
      RECT 604.1000 660.1450 609.2500 663.1450 ;
      RECT 595.9500 660.1450 601.1000 663.1450 ;
      RECT 587.8000 660.1450 592.9500 663.1450 ;
      RECT 579.6500 660.1450 584.8000 663.1450 ;
      RECT 571.5000 660.1450 576.6500 663.1450 ;
      RECT 563.3500 660.1450 568.5000 663.1450 ;
      RECT 555.2000 660.1450 560.3500 663.1450 ;
      RECT 547.0500 660.1450 552.2000 663.1450 ;
      RECT 538.9000 660.1450 544.0500 663.1450 ;
      RECT 530.7500 660.1450 535.9000 663.1450 ;
      RECT 522.6000 660.1450 527.7500 663.1450 ;
      RECT 514.4500 660.1450 519.6000 663.1450 ;
      RECT 506.3000 660.1450 511.4500 663.1450 ;
      RECT 498.1500 660.1450 503.3000 663.1450 ;
      RECT 490.0000 660.1450 495.1500 663.1450 ;
      RECT 481.8500 660.1450 487.0000 663.1450 ;
      RECT 473.7000 660.1450 478.8500 663.1450 ;
      RECT 465.5500 660.1450 470.7000 663.1450 ;
      RECT 457.4000 660.1450 462.5500 663.1450 ;
      RECT 449.2500 660.1450 454.4000 663.1450 ;
      RECT 441.1000 660.1450 446.2500 663.1450 ;
      RECT 432.9500 660.1450 438.1000 663.1450 ;
      RECT 424.8000 660.1450 429.9500 663.1450 ;
      RECT 416.6500 660.1450 421.8000 663.1450 ;
      RECT 396.5000 660.1450 413.6500 663.1450 ;
      RECT 346.5000 660.1450 393.5000 663.1450 ;
      RECT 326.4650 660.1450 343.5000 663.1450 ;
      RECT 317.9500 660.1450 323.4650 663.1450 ;
      RECT 309.4350 660.1450 314.9500 663.1450 ;
      RECT 300.9200 660.1450 306.4350 663.1450 ;
      RECT 292.4050 660.1450 297.9200 663.1450 ;
      RECT 283.8900 660.1450 289.4050 663.1450 ;
      RECT 275.3750 660.1450 280.8900 663.1450 ;
      RECT 266.8600 660.1450 272.3750 663.1450 ;
      RECT 258.3450 660.1450 263.8600 663.1450 ;
      RECT 249.8300 660.1450 255.3450 663.1450 ;
      RECT 241.3150 660.1450 246.8300 663.1450 ;
      RECT 232.8000 660.1450 238.3150 663.1450 ;
      RECT 224.2850 660.1450 229.8000 663.1450 ;
      RECT 215.7700 660.1450 221.2850 663.1450 ;
      RECT 207.2550 660.1450 212.7700 663.1450 ;
      RECT 198.7400 660.1450 204.2550 663.1450 ;
      RECT 190.2250 660.1450 195.7400 663.1450 ;
      RECT 181.7100 660.1450 187.2250 663.1450 ;
      RECT 173.1950 660.1450 178.7100 663.1450 ;
      RECT 164.6800 660.1450 170.1950 663.1450 ;
      RECT 156.1650 660.1450 161.6800 663.1450 ;
      RECT 147.6500 660.1450 153.1650 663.1450 ;
      RECT 139.1350 660.1450 144.6500 663.1450 ;
      RECT 130.6200 660.1450 136.1350 663.1450 ;
      RECT 122.1050 660.1450 127.6200 663.1450 ;
      RECT 113.5900 660.1450 119.1050 663.1450 ;
      RECT 105.0750 660.1450 110.5900 663.1450 ;
      RECT 96.5600 660.1450 102.0750 663.1450 ;
      RECT 88.0450 660.1450 93.5600 663.1450 ;
      RECT 79.5300 660.1450 85.0450 663.1450 ;
      RECT 71.0150 660.1450 76.5300 663.1450 ;
      RECT 62.5000 660.1450 68.0150 663.1450 ;
      RECT 46.5000 660.1450 59.5000 663.1450 ;
      RECT 8.5000 660.1450 43.5000 663.1450 ;
      RECT 0.0000 660.1450 5.5000 663.1450 ;
      RECT 0.0000 658.7000 1120.0000 660.1450 ;
      RECT 1116.6000 658.1450 1120.0000 658.7000 ;
      RECT 0.0000 656.0500 1113.6000 658.7000 ;
      RECT 1118.5000 655.1450 1120.0000 658.1450 ;
      RECT 1114.5000 653.0500 1120.0000 655.1450 ;
      RECT 1076.5000 653.0500 1111.5000 656.0500 ;
      RECT 1060.5000 653.0500 1073.5000 656.0500 ;
      RECT 1052.3500 653.0500 1057.5000 656.0500 ;
      RECT 1044.2000 653.0500 1049.3500 656.0500 ;
      RECT 1036.0500 653.0500 1041.2000 656.0500 ;
      RECT 1027.9000 653.0500 1033.0500 656.0500 ;
      RECT 1019.7500 653.0500 1024.9000 656.0500 ;
      RECT 1011.6000 653.0500 1016.7500 656.0500 ;
      RECT 1003.4500 653.0500 1008.6000 656.0500 ;
      RECT 995.3000 653.0500 1000.4500 656.0500 ;
      RECT 987.1500 653.0500 992.3000 656.0500 ;
      RECT 979.0000 653.0500 984.1500 656.0500 ;
      RECT 970.8500 653.0500 976.0000 656.0500 ;
      RECT 962.7000 653.0500 967.8500 656.0500 ;
      RECT 954.5500 653.0500 959.7000 656.0500 ;
      RECT 946.4000 653.0500 951.5500 656.0500 ;
      RECT 938.2500 653.0500 943.4000 656.0500 ;
      RECT 930.1000 653.0500 935.2500 656.0500 ;
      RECT 921.9500 653.0500 927.1000 656.0500 ;
      RECT 913.8000 653.0500 918.9500 656.0500 ;
      RECT 905.6500 653.0500 910.8000 656.0500 ;
      RECT 897.5000 653.0500 902.6500 656.0500 ;
      RECT 889.3500 653.0500 894.5000 656.0500 ;
      RECT 881.2000 653.0500 886.3500 656.0500 ;
      RECT 873.0500 653.0500 878.2000 656.0500 ;
      RECT 864.9000 653.0500 870.0500 656.0500 ;
      RECT 856.7500 653.0500 861.9000 656.0500 ;
      RECT 848.6000 653.0500 853.7500 656.0500 ;
      RECT 840.4500 653.0500 845.6000 656.0500 ;
      RECT 832.3000 653.0500 837.4500 656.0500 ;
      RECT 824.1500 653.0500 829.3000 656.0500 ;
      RECT 816.0000 653.0500 821.1500 656.0500 ;
      RECT 807.8500 653.0500 813.0000 656.0500 ;
      RECT 799.7000 653.0500 804.8500 656.0500 ;
      RECT 791.5500 653.0500 796.7000 656.0500 ;
      RECT 783.4000 653.0500 788.5500 656.0500 ;
      RECT 775.2500 653.0500 780.4000 656.0500 ;
      RECT 767.1000 653.0500 772.2500 656.0500 ;
      RECT 758.9500 653.0500 764.1000 656.0500 ;
      RECT 750.8000 653.0500 755.9500 656.0500 ;
      RECT 742.6500 653.0500 747.8000 656.0500 ;
      RECT 734.5000 653.0500 739.6500 656.0500 ;
      RECT 726.3500 653.0500 731.5000 656.0500 ;
      RECT 718.2000 653.0500 723.3500 656.0500 ;
      RECT 710.0500 653.0500 715.2000 656.0500 ;
      RECT 701.9000 653.0500 707.0500 656.0500 ;
      RECT 693.7500 653.0500 698.9000 656.0500 ;
      RECT 685.6000 653.0500 690.7500 656.0500 ;
      RECT 677.4500 653.0500 682.6000 656.0500 ;
      RECT 669.3000 653.0500 674.4500 656.0500 ;
      RECT 661.1500 653.0500 666.3000 656.0500 ;
      RECT 653.0000 653.0500 658.1500 656.0500 ;
      RECT 644.8500 653.0500 650.0000 656.0500 ;
      RECT 636.7000 653.0500 641.8500 656.0500 ;
      RECT 628.5500 653.0500 633.7000 656.0500 ;
      RECT 620.4000 653.0500 625.5500 656.0500 ;
      RECT 612.2500 653.0500 617.4000 656.0500 ;
      RECT 604.1000 653.0500 609.2500 656.0500 ;
      RECT 595.9500 653.0500 601.1000 656.0500 ;
      RECT 587.8000 653.0500 592.9500 656.0500 ;
      RECT 579.6500 653.0500 584.8000 656.0500 ;
      RECT 571.5000 653.0500 576.6500 656.0500 ;
      RECT 563.3500 653.0500 568.5000 656.0500 ;
      RECT 555.2000 653.0500 560.3500 656.0500 ;
      RECT 547.0500 653.0500 552.2000 656.0500 ;
      RECT 538.9000 653.0500 544.0500 656.0500 ;
      RECT 530.7500 653.0500 535.9000 656.0500 ;
      RECT 522.6000 653.0500 527.7500 656.0500 ;
      RECT 514.4500 653.0500 519.6000 656.0500 ;
      RECT 506.3000 653.0500 511.4500 656.0500 ;
      RECT 498.1500 653.0500 503.3000 656.0500 ;
      RECT 490.0000 653.0500 495.1500 656.0500 ;
      RECT 481.8500 653.0500 487.0000 656.0500 ;
      RECT 473.7000 653.0500 478.8500 656.0500 ;
      RECT 465.5500 653.0500 470.7000 656.0500 ;
      RECT 457.4000 653.0500 462.5500 656.0500 ;
      RECT 449.2500 653.0500 454.4000 656.0500 ;
      RECT 441.1000 653.0500 446.2500 656.0500 ;
      RECT 432.9500 653.0500 438.1000 656.0500 ;
      RECT 424.8000 653.0500 429.9500 656.0500 ;
      RECT 416.6500 653.0500 421.8000 656.0500 ;
      RECT 396.5000 653.0500 413.6500 656.0500 ;
      RECT 346.5000 653.0500 393.5000 656.0500 ;
      RECT 326.4650 653.0500 343.5000 656.0500 ;
      RECT 317.9500 653.0500 323.4650 656.0500 ;
      RECT 309.4350 653.0500 314.9500 656.0500 ;
      RECT 300.9200 653.0500 306.4350 656.0500 ;
      RECT 292.4050 653.0500 297.9200 656.0500 ;
      RECT 283.8900 653.0500 289.4050 656.0500 ;
      RECT 275.3750 653.0500 280.8900 656.0500 ;
      RECT 266.8600 653.0500 272.3750 656.0500 ;
      RECT 258.3450 653.0500 263.8600 656.0500 ;
      RECT 249.8300 653.0500 255.3450 656.0500 ;
      RECT 241.3150 653.0500 246.8300 656.0500 ;
      RECT 232.8000 653.0500 238.3150 656.0500 ;
      RECT 224.2850 653.0500 229.8000 656.0500 ;
      RECT 215.7700 653.0500 221.2850 656.0500 ;
      RECT 207.2550 653.0500 212.7700 656.0500 ;
      RECT 198.7400 653.0500 204.2550 656.0500 ;
      RECT 190.2250 653.0500 195.7400 656.0500 ;
      RECT 181.7100 653.0500 187.2250 656.0500 ;
      RECT 173.1950 653.0500 178.7100 656.0500 ;
      RECT 164.6800 653.0500 170.1950 656.0500 ;
      RECT 156.1650 653.0500 161.6800 656.0500 ;
      RECT 147.6500 653.0500 153.1650 656.0500 ;
      RECT 139.1350 653.0500 144.6500 656.0500 ;
      RECT 130.6200 653.0500 136.1350 656.0500 ;
      RECT 122.1050 653.0500 127.6200 656.0500 ;
      RECT 113.5900 653.0500 119.1050 656.0500 ;
      RECT 105.0750 653.0500 110.5900 656.0500 ;
      RECT 96.5600 653.0500 102.0750 656.0500 ;
      RECT 88.0450 653.0500 93.5600 656.0500 ;
      RECT 79.5300 653.0500 85.0450 656.0500 ;
      RECT 71.0150 653.0500 76.5300 656.0500 ;
      RECT 62.5000 653.0500 68.0150 656.0500 ;
      RECT 46.5000 653.0500 59.5000 656.0500 ;
      RECT 8.5000 653.0500 43.5000 656.0500 ;
      RECT 0.0000 653.0500 5.5000 656.0500 ;
      RECT 0.0000 651.5000 1120.0000 653.0500 ;
      RECT 1116.6000 651.0500 1120.0000 651.5000 ;
      RECT 0.0000 648.9550 1113.6000 651.5000 ;
      RECT 1118.5000 648.0500 1120.0000 651.0500 ;
      RECT 1114.5000 645.9550 1120.0000 648.0500 ;
      RECT 1076.5000 645.9550 1111.5000 648.9550 ;
      RECT 1060.5000 645.9550 1073.5000 648.9550 ;
      RECT 1052.3500 645.9550 1057.5000 648.9550 ;
      RECT 1044.2000 645.9550 1049.3500 648.9550 ;
      RECT 1036.0500 645.9550 1041.2000 648.9550 ;
      RECT 1027.9000 645.9550 1033.0500 648.9550 ;
      RECT 1019.7500 645.9550 1024.9000 648.9550 ;
      RECT 1011.6000 645.9550 1016.7500 648.9550 ;
      RECT 1003.4500 645.9550 1008.6000 648.9550 ;
      RECT 995.3000 645.9550 1000.4500 648.9550 ;
      RECT 987.1500 645.9550 992.3000 648.9550 ;
      RECT 979.0000 645.9550 984.1500 648.9550 ;
      RECT 970.8500 645.9550 976.0000 648.9550 ;
      RECT 962.7000 645.9550 967.8500 648.9550 ;
      RECT 954.5500 645.9550 959.7000 648.9550 ;
      RECT 946.4000 645.9550 951.5500 648.9550 ;
      RECT 938.2500 645.9550 943.4000 648.9550 ;
      RECT 930.1000 645.9550 935.2500 648.9550 ;
      RECT 921.9500 645.9550 927.1000 648.9550 ;
      RECT 913.8000 645.9550 918.9500 648.9550 ;
      RECT 905.6500 645.9550 910.8000 648.9550 ;
      RECT 897.5000 645.9550 902.6500 648.9550 ;
      RECT 889.3500 645.9550 894.5000 648.9550 ;
      RECT 881.2000 645.9550 886.3500 648.9550 ;
      RECT 873.0500 645.9550 878.2000 648.9550 ;
      RECT 864.9000 645.9550 870.0500 648.9550 ;
      RECT 856.7500 645.9550 861.9000 648.9550 ;
      RECT 848.6000 645.9550 853.7500 648.9550 ;
      RECT 840.4500 645.9550 845.6000 648.9550 ;
      RECT 832.3000 645.9550 837.4500 648.9550 ;
      RECT 824.1500 645.9550 829.3000 648.9550 ;
      RECT 816.0000 645.9550 821.1500 648.9550 ;
      RECT 807.8500 645.9550 813.0000 648.9550 ;
      RECT 799.7000 645.9550 804.8500 648.9550 ;
      RECT 791.5500 645.9550 796.7000 648.9550 ;
      RECT 783.4000 645.9550 788.5500 648.9550 ;
      RECT 775.2500 645.9550 780.4000 648.9550 ;
      RECT 767.1000 645.9550 772.2500 648.9550 ;
      RECT 758.9500 645.9550 764.1000 648.9550 ;
      RECT 750.8000 645.9550 755.9500 648.9550 ;
      RECT 742.6500 645.9550 747.8000 648.9550 ;
      RECT 734.5000 645.9550 739.6500 648.9550 ;
      RECT 726.3500 645.9550 731.5000 648.9550 ;
      RECT 718.2000 645.9550 723.3500 648.9550 ;
      RECT 710.0500 645.9550 715.2000 648.9550 ;
      RECT 701.9000 645.9550 707.0500 648.9550 ;
      RECT 693.7500 645.9550 698.9000 648.9550 ;
      RECT 685.6000 645.9550 690.7500 648.9550 ;
      RECT 677.4500 645.9550 682.6000 648.9550 ;
      RECT 669.3000 645.9550 674.4500 648.9550 ;
      RECT 661.1500 645.9550 666.3000 648.9550 ;
      RECT 653.0000 645.9550 658.1500 648.9550 ;
      RECT 644.8500 645.9550 650.0000 648.9550 ;
      RECT 636.7000 645.9550 641.8500 648.9550 ;
      RECT 628.5500 645.9550 633.7000 648.9550 ;
      RECT 620.4000 645.9550 625.5500 648.9550 ;
      RECT 612.2500 645.9550 617.4000 648.9550 ;
      RECT 604.1000 645.9550 609.2500 648.9550 ;
      RECT 595.9500 645.9550 601.1000 648.9550 ;
      RECT 587.8000 645.9550 592.9500 648.9550 ;
      RECT 579.6500 645.9550 584.8000 648.9550 ;
      RECT 571.5000 645.9550 576.6500 648.9550 ;
      RECT 563.3500 645.9550 568.5000 648.9550 ;
      RECT 555.2000 645.9550 560.3500 648.9550 ;
      RECT 547.0500 645.9550 552.2000 648.9550 ;
      RECT 538.9000 645.9550 544.0500 648.9550 ;
      RECT 530.7500 645.9550 535.9000 648.9550 ;
      RECT 522.6000 645.9550 527.7500 648.9550 ;
      RECT 514.4500 645.9550 519.6000 648.9550 ;
      RECT 506.3000 645.9550 511.4500 648.9550 ;
      RECT 498.1500 645.9550 503.3000 648.9550 ;
      RECT 490.0000 645.9550 495.1500 648.9550 ;
      RECT 481.8500 645.9550 487.0000 648.9550 ;
      RECT 473.7000 645.9550 478.8500 648.9550 ;
      RECT 465.5500 645.9550 470.7000 648.9550 ;
      RECT 457.4000 645.9550 462.5500 648.9550 ;
      RECT 449.2500 645.9550 454.4000 648.9550 ;
      RECT 441.1000 645.9550 446.2500 648.9550 ;
      RECT 432.9500 645.9550 438.1000 648.9550 ;
      RECT 424.8000 645.9550 429.9500 648.9550 ;
      RECT 416.6500 645.9550 421.8000 648.9550 ;
      RECT 396.5000 645.9550 413.6500 648.9550 ;
      RECT 346.5000 645.9550 393.5000 648.9550 ;
      RECT 326.4650 645.9550 343.5000 648.9550 ;
      RECT 317.9500 645.9550 323.4650 648.9550 ;
      RECT 309.4350 645.9550 314.9500 648.9550 ;
      RECT 300.9200 645.9550 306.4350 648.9550 ;
      RECT 292.4050 645.9550 297.9200 648.9550 ;
      RECT 283.8900 645.9550 289.4050 648.9550 ;
      RECT 275.3750 645.9550 280.8900 648.9550 ;
      RECT 266.8600 645.9550 272.3750 648.9550 ;
      RECT 258.3450 645.9550 263.8600 648.9550 ;
      RECT 249.8300 645.9550 255.3450 648.9550 ;
      RECT 241.3150 645.9550 246.8300 648.9550 ;
      RECT 232.8000 645.9550 238.3150 648.9550 ;
      RECT 224.2850 645.9550 229.8000 648.9550 ;
      RECT 215.7700 645.9550 221.2850 648.9550 ;
      RECT 207.2550 645.9550 212.7700 648.9550 ;
      RECT 198.7400 645.9550 204.2550 648.9550 ;
      RECT 190.2250 645.9550 195.7400 648.9550 ;
      RECT 181.7100 645.9550 187.2250 648.9550 ;
      RECT 173.1950 645.9550 178.7100 648.9550 ;
      RECT 164.6800 645.9550 170.1950 648.9550 ;
      RECT 156.1650 645.9550 161.6800 648.9550 ;
      RECT 147.6500 645.9550 153.1650 648.9550 ;
      RECT 139.1350 645.9550 144.6500 648.9550 ;
      RECT 130.6200 645.9550 136.1350 648.9550 ;
      RECT 122.1050 645.9550 127.6200 648.9550 ;
      RECT 113.5900 645.9550 119.1050 648.9550 ;
      RECT 105.0750 645.9550 110.5900 648.9550 ;
      RECT 96.5600 645.9550 102.0750 648.9550 ;
      RECT 88.0450 645.9550 93.5600 648.9550 ;
      RECT 79.5300 645.9550 85.0450 648.9550 ;
      RECT 71.0150 645.9550 76.5300 648.9550 ;
      RECT 62.5000 645.9550 68.0150 648.9550 ;
      RECT 46.5000 645.9550 59.5000 648.9550 ;
      RECT 8.5000 645.9550 43.5000 648.9550 ;
      RECT 0.0000 645.9550 5.5000 648.9550 ;
      RECT 0.0000 644.5000 1120.0000 645.9550 ;
      RECT 1116.6000 643.9550 1120.0000 644.5000 ;
      RECT 0.0000 641.8600 1113.6000 644.5000 ;
      RECT 1118.5000 640.9550 1120.0000 643.9550 ;
      RECT 1114.5000 638.8600 1120.0000 640.9550 ;
      RECT 1076.5000 638.8600 1111.5000 641.8600 ;
      RECT 1060.5000 638.8600 1073.5000 641.8600 ;
      RECT 1052.3500 638.8600 1057.5000 641.8600 ;
      RECT 1044.2000 638.8600 1049.3500 641.8600 ;
      RECT 1036.0500 638.8600 1041.2000 641.8600 ;
      RECT 1027.9000 638.8600 1033.0500 641.8600 ;
      RECT 1019.7500 638.8600 1024.9000 641.8600 ;
      RECT 1011.6000 638.8600 1016.7500 641.8600 ;
      RECT 1003.4500 638.8600 1008.6000 641.8600 ;
      RECT 995.3000 638.8600 1000.4500 641.8600 ;
      RECT 987.1500 638.8600 992.3000 641.8600 ;
      RECT 979.0000 638.8600 984.1500 641.8600 ;
      RECT 970.8500 638.8600 976.0000 641.8600 ;
      RECT 962.7000 638.8600 967.8500 641.8600 ;
      RECT 954.5500 638.8600 959.7000 641.8600 ;
      RECT 946.4000 638.8600 951.5500 641.8600 ;
      RECT 938.2500 638.8600 943.4000 641.8600 ;
      RECT 930.1000 638.8600 935.2500 641.8600 ;
      RECT 921.9500 638.8600 927.1000 641.8600 ;
      RECT 913.8000 638.8600 918.9500 641.8600 ;
      RECT 905.6500 638.8600 910.8000 641.8600 ;
      RECT 897.5000 638.8600 902.6500 641.8600 ;
      RECT 889.3500 638.8600 894.5000 641.8600 ;
      RECT 881.2000 638.8600 886.3500 641.8600 ;
      RECT 873.0500 638.8600 878.2000 641.8600 ;
      RECT 864.9000 638.8600 870.0500 641.8600 ;
      RECT 856.7500 638.8600 861.9000 641.8600 ;
      RECT 848.6000 638.8600 853.7500 641.8600 ;
      RECT 840.4500 638.8600 845.6000 641.8600 ;
      RECT 832.3000 638.8600 837.4500 641.8600 ;
      RECT 824.1500 638.8600 829.3000 641.8600 ;
      RECT 816.0000 638.8600 821.1500 641.8600 ;
      RECT 807.8500 638.8600 813.0000 641.8600 ;
      RECT 799.7000 638.8600 804.8500 641.8600 ;
      RECT 791.5500 638.8600 796.7000 641.8600 ;
      RECT 783.4000 638.8600 788.5500 641.8600 ;
      RECT 775.2500 638.8600 780.4000 641.8600 ;
      RECT 767.1000 638.8600 772.2500 641.8600 ;
      RECT 758.9500 638.8600 764.1000 641.8600 ;
      RECT 750.8000 638.8600 755.9500 641.8600 ;
      RECT 742.6500 638.8600 747.8000 641.8600 ;
      RECT 734.5000 638.8600 739.6500 641.8600 ;
      RECT 726.3500 638.8600 731.5000 641.8600 ;
      RECT 718.2000 638.8600 723.3500 641.8600 ;
      RECT 710.0500 638.8600 715.2000 641.8600 ;
      RECT 701.9000 638.8600 707.0500 641.8600 ;
      RECT 693.7500 638.8600 698.9000 641.8600 ;
      RECT 685.6000 638.8600 690.7500 641.8600 ;
      RECT 677.4500 638.8600 682.6000 641.8600 ;
      RECT 669.3000 638.8600 674.4500 641.8600 ;
      RECT 661.1500 638.8600 666.3000 641.8600 ;
      RECT 653.0000 638.8600 658.1500 641.8600 ;
      RECT 644.8500 638.8600 650.0000 641.8600 ;
      RECT 636.7000 638.8600 641.8500 641.8600 ;
      RECT 628.5500 638.8600 633.7000 641.8600 ;
      RECT 620.4000 638.8600 625.5500 641.8600 ;
      RECT 612.2500 638.8600 617.4000 641.8600 ;
      RECT 604.1000 638.8600 609.2500 641.8600 ;
      RECT 595.9500 638.8600 601.1000 641.8600 ;
      RECT 587.8000 638.8600 592.9500 641.8600 ;
      RECT 579.6500 638.8600 584.8000 641.8600 ;
      RECT 571.5000 638.8600 576.6500 641.8600 ;
      RECT 563.3500 638.8600 568.5000 641.8600 ;
      RECT 555.2000 638.8600 560.3500 641.8600 ;
      RECT 547.0500 638.8600 552.2000 641.8600 ;
      RECT 538.9000 638.8600 544.0500 641.8600 ;
      RECT 530.7500 638.8600 535.9000 641.8600 ;
      RECT 522.6000 638.8600 527.7500 641.8600 ;
      RECT 514.4500 638.8600 519.6000 641.8600 ;
      RECT 506.3000 638.8600 511.4500 641.8600 ;
      RECT 498.1500 638.8600 503.3000 641.8600 ;
      RECT 490.0000 638.8600 495.1500 641.8600 ;
      RECT 481.8500 638.8600 487.0000 641.8600 ;
      RECT 473.7000 638.8600 478.8500 641.8600 ;
      RECT 465.5500 638.8600 470.7000 641.8600 ;
      RECT 457.4000 638.8600 462.5500 641.8600 ;
      RECT 449.2500 638.8600 454.4000 641.8600 ;
      RECT 441.1000 638.8600 446.2500 641.8600 ;
      RECT 432.9500 638.8600 438.1000 641.8600 ;
      RECT 424.8000 638.8600 429.9500 641.8600 ;
      RECT 416.6500 638.8600 421.8000 641.8600 ;
      RECT 396.5000 638.8600 413.6500 641.8600 ;
      RECT 346.5000 638.8600 393.5000 641.8600 ;
      RECT 326.4650 638.8600 343.5000 641.8600 ;
      RECT 317.9500 638.8600 323.4650 641.8600 ;
      RECT 309.4350 638.8600 314.9500 641.8600 ;
      RECT 300.9200 638.8600 306.4350 641.8600 ;
      RECT 292.4050 638.8600 297.9200 641.8600 ;
      RECT 283.8900 638.8600 289.4050 641.8600 ;
      RECT 275.3750 638.8600 280.8900 641.8600 ;
      RECT 266.8600 638.8600 272.3750 641.8600 ;
      RECT 258.3450 638.8600 263.8600 641.8600 ;
      RECT 249.8300 638.8600 255.3450 641.8600 ;
      RECT 241.3150 638.8600 246.8300 641.8600 ;
      RECT 232.8000 638.8600 238.3150 641.8600 ;
      RECT 224.2850 638.8600 229.8000 641.8600 ;
      RECT 215.7700 638.8600 221.2850 641.8600 ;
      RECT 207.2550 638.8600 212.7700 641.8600 ;
      RECT 198.7400 638.8600 204.2550 641.8600 ;
      RECT 190.2250 638.8600 195.7400 641.8600 ;
      RECT 181.7100 638.8600 187.2250 641.8600 ;
      RECT 173.1950 638.8600 178.7100 641.8600 ;
      RECT 164.6800 638.8600 170.1950 641.8600 ;
      RECT 156.1650 638.8600 161.6800 641.8600 ;
      RECT 147.6500 638.8600 153.1650 641.8600 ;
      RECT 139.1350 638.8600 144.6500 641.8600 ;
      RECT 130.6200 638.8600 136.1350 641.8600 ;
      RECT 122.1050 638.8600 127.6200 641.8600 ;
      RECT 113.5900 638.8600 119.1050 641.8600 ;
      RECT 105.0750 638.8600 110.5900 641.8600 ;
      RECT 96.5600 638.8600 102.0750 641.8600 ;
      RECT 88.0450 638.8600 93.5600 641.8600 ;
      RECT 79.5300 638.8600 85.0450 641.8600 ;
      RECT 71.0150 638.8600 76.5300 641.8600 ;
      RECT 62.5000 638.8600 68.0150 641.8600 ;
      RECT 46.5000 638.8600 59.5000 641.8600 ;
      RECT 8.5000 638.8600 43.5000 641.8600 ;
      RECT 0.0000 638.8600 5.5000 641.8600 ;
      RECT 0.0000 637.3000 1120.0000 638.8600 ;
      RECT 1116.6000 636.8600 1120.0000 637.3000 ;
      RECT 0.0000 634.7650 1113.6000 637.3000 ;
      RECT 1118.5000 633.8600 1120.0000 636.8600 ;
      RECT 1114.5000 631.7650 1120.0000 633.8600 ;
      RECT 1076.5000 631.7650 1111.5000 634.7650 ;
      RECT 1060.5000 631.7650 1073.5000 634.7650 ;
      RECT 1052.3500 631.7650 1057.5000 634.7650 ;
      RECT 1044.2000 631.7650 1049.3500 634.7650 ;
      RECT 1036.0500 631.7650 1041.2000 634.7650 ;
      RECT 1027.9000 631.7650 1033.0500 634.7650 ;
      RECT 1019.7500 631.7650 1024.9000 634.7650 ;
      RECT 1011.6000 631.7650 1016.7500 634.7650 ;
      RECT 1003.4500 631.7650 1008.6000 634.7650 ;
      RECT 995.3000 631.7650 1000.4500 634.7650 ;
      RECT 987.1500 631.7650 992.3000 634.7650 ;
      RECT 979.0000 631.7650 984.1500 634.7650 ;
      RECT 970.8500 631.7650 976.0000 634.7650 ;
      RECT 962.7000 631.7650 967.8500 634.7650 ;
      RECT 954.5500 631.7650 959.7000 634.7650 ;
      RECT 946.4000 631.7650 951.5500 634.7650 ;
      RECT 938.2500 631.7650 943.4000 634.7650 ;
      RECT 930.1000 631.7650 935.2500 634.7650 ;
      RECT 921.9500 631.7650 927.1000 634.7650 ;
      RECT 913.8000 631.7650 918.9500 634.7650 ;
      RECT 905.6500 631.7650 910.8000 634.7650 ;
      RECT 897.5000 631.7650 902.6500 634.7650 ;
      RECT 889.3500 631.7650 894.5000 634.7650 ;
      RECT 881.2000 631.7650 886.3500 634.7650 ;
      RECT 873.0500 631.7650 878.2000 634.7650 ;
      RECT 864.9000 631.7650 870.0500 634.7650 ;
      RECT 856.7500 631.7650 861.9000 634.7650 ;
      RECT 848.6000 631.7650 853.7500 634.7650 ;
      RECT 840.4500 631.7650 845.6000 634.7650 ;
      RECT 832.3000 631.7650 837.4500 634.7650 ;
      RECT 824.1500 631.7650 829.3000 634.7650 ;
      RECT 816.0000 631.7650 821.1500 634.7650 ;
      RECT 807.8500 631.7650 813.0000 634.7650 ;
      RECT 799.7000 631.7650 804.8500 634.7650 ;
      RECT 791.5500 631.7650 796.7000 634.7650 ;
      RECT 783.4000 631.7650 788.5500 634.7650 ;
      RECT 775.2500 631.7650 780.4000 634.7650 ;
      RECT 767.1000 631.7650 772.2500 634.7650 ;
      RECT 758.9500 631.7650 764.1000 634.7650 ;
      RECT 750.8000 631.7650 755.9500 634.7650 ;
      RECT 742.6500 631.7650 747.8000 634.7650 ;
      RECT 734.5000 631.7650 739.6500 634.7650 ;
      RECT 726.3500 631.7650 731.5000 634.7650 ;
      RECT 718.2000 631.7650 723.3500 634.7650 ;
      RECT 710.0500 631.7650 715.2000 634.7650 ;
      RECT 701.9000 631.7650 707.0500 634.7650 ;
      RECT 693.7500 631.7650 698.9000 634.7650 ;
      RECT 685.6000 631.7650 690.7500 634.7650 ;
      RECT 677.4500 631.7650 682.6000 634.7650 ;
      RECT 669.3000 631.7650 674.4500 634.7650 ;
      RECT 661.1500 631.7650 666.3000 634.7650 ;
      RECT 653.0000 631.7650 658.1500 634.7650 ;
      RECT 644.8500 631.7650 650.0000 634.7650 ;
      RECT 636.7000 631.7650 641.8500 634.7650 ;
      RECT 628.5500 631.7650 633.7000 634.7650 ;
      RECT 620.4000 631.7650 625.5500 634.7650 ;
      RECT 612.2500 631.7650 617.4000 634.7650 ;
      RECT 604.1000 631.7650 609.2500 634.7650 ;
      RECT 595.9500 631.7650 601.1000 634.7650 ;
      RECT 587.8000 631.7650 592.9500 634.7650 ;
      RECT 579.6500 631.7650 584.8000 634.7650 ;
      RECT 571.5000 631.7650 576.6500 634.7650 ;
      RECT 563.3500 631.7650 568.5000 634.7650 ;
      RECT 555.2000 631.7650 560.3500 634.7650 ;
      RECT 547.0500 631.7650 552.2000 634.7650 ;
      RECT 538.9000 631.7650 544.0500 634.7650 ;
      RECT 530.7500 631.7650 535.9000 634.7650 ;
      RECT 522.6000 631.7650 527.7500 634.7650 ;
      RECT 514.4500 631.7650 519.6000 634.7650 ;
      RECT 506.3000 631.7650 511.4500 634.7650 ;
      RECT 498.1500 631.7650 503.3000 634.7650 ;
      RECT 490.0000 631.7650 495.1500 634.7650 ;
      RECT 481.8500 631.7650 487.0000 634.7650 ;
      RECT 473.7000 631.7650 478.8500 634.7650 ;
      RECT 465.5500 631.7650 470.7000 634.7650 ;
      RECT 457.4000 631.7650 462.5500 634.7650 ;
      RECT 449.2500 631.7650 454.4000 634.7650 ;
      RECT 441.1000 631.7650 446.2500 634.7650 ;
      RECT 432.9500 631.7650 438.1000 634.7650 ;
      RECT 424.8000 631.7650 429.9500 634.7650 ;
      RECT 416.6500 631.7650 421.8000 634.7650 ;
      RECT 396.5000 631.7650 413.6500 634.7650 ;
      RECT 346.5000 631.7650 393.5000 634.7650 ;
      RECT 326.4650 631.7650 343.5000 634.7650 ;
      RECT 317.9500 631.7650 323.4650 634.7650 ;
      RECT 309.4350 631.7650 314.9500 634.7650 ;
      RECT 300.9200 631.7650 306.4350 634.7650 ;
      RECT 292.4050 631.7650 297.9200 634.7650 ;
      RECT 283.8900 631.7650 289.4050 634.7650 ;
      RECT 275.3750 631.7650 280.8900 634.7650 ;
      RECT 266.8600 631.7650 272.3750 634.7650 ;
      RECT 258.3450 631.7650 263.8600 634.7650 ;
      RECT 249.8300 631.7650 255.3450 634.7650 ;
      RECT 241.3150 631.7650 246.8300 634.7650 ;
      RECT 232.8000 631.7650 238.3150 634.7650 ;
      RECT 224.2850 631.7650 229.8000 634.7650 ;
      RECT 215.7700 631.7650 221.2850 634.7650 ;
      RECT 207.2550 631.7650 212.7700 634.7650 ;
      RECT 198.7400 631.7650 204.2550 634.7650 ;
      RECT 190.2250 631.7650 195.7400 634.7650 ;
      RECT 181.7100 631.7650 187.2250 634.7650 ;
      RECT 173.1950 631.7650 178.7100 634.7650 ;
      RECT 164.6800 631.7650 170.1950 634.7650 ;
      RECT 156.1650 631.7650 161.6800 634.7650 ;
      RECT 147.6500 631.7650 153.1650 634.7650 ;
      RECT 139.1350 631.7650 144.6500 634.7650 ;
      RECT 130.6200 631.7650 136.1350 634.7650 ;
      RECT 122.1050 631.7650 127.6200 634.7650 ;
      RECT 113.5900 631.7650 119.1050 634.7650 ;
      RECT 105.0750 631.7650 110.5900 634.7650 ;
      RECT 96.5600 631.7650 102.0750 634.7650 ;
      RECT 88.0450 631.7650 93.5600 634.7650 ;
      RECT 79.5300 631.7650 85.0450 634.7650 ;
      RECT 71.0150 631.7650 76.5300 634.7650 ;
      RECT 62.5000 631.7650 68.0150 634.7650 ;
      RECT 46.5000 631.7650 59.5000 634.7650 ;
      RECT 8.5000 631.7650 43.5000 634.7650 ;
      RECT 0.0000 631.7650 5.5000 634.7650 ;
      RECT 0.0000 630.3000 1120.0000 631.7650 ;
      RECT 1116.6000 629.7650 1120.0000 630.3000 ;
      RECT 0.0000 627.6700 1113.6000 630.3000 ;
      RECT 1118.5000 626.7650 1120.0000 629.7650 ;
      RECT 1114.5000 624.6700 1120.0000 626.7650 ;
      RECT 1076.5000 624.6700 1111.5000 627.6700 ;
      RECT 1060.5000 624.6700 1073.5000 627.6700 ;
      RECT 1052.3500 624.6700 1057.5000 627.6700 ;
      RECT 1044.2000 624.6700 1049.3500 627.6700 ;
      RECT 1036.0500 624.6700 1041.2000 627.6700 ;
      RECT 1027.9000 624.6700 1033.0500 627.6700 ;
      RECT 1019.7500 624.6700 1024.9000 627.6700 ;
      RECT 1011.6000 624.6700 1016.7500 627.6700 ;
      RECT 1003.4500 624.6700 1008.6000 627.6700 ;
      RECT 995.3000 624.6700 1000.4500 627.6700 ;
      RECT 987.1500 624.6700 992.3000 627.6700 ;
      RECT 979.0000 624.6700 984.1500 627.6700 ;
      RECT 970.8500 624.6700 976.0000 627.6700 ;
      RECT 962.7000 624.6700 967.8500 627.6700 ;
      RECT 954.5500 624.6700 959.7000 627.6700 ;
      RECT 946.4000 624.6700 951.5500 627.6700 ;
      RECT 938.2500 624.6700 943.4000 627.6700 ;
      RECT 930.1000 624.6700 935.2500 627.6700 ;
      RECT 921.9500 624.6700 927.1000 627.6700 ;
      RECT 913.8000 624.6700 918.9500 627.6700 ;
      RECT 905.6500 624.6700 910.8000 627.6700 ;
      RECT 897.5000 624.6700 902.6500 627.6700 ;
      RECT 889.3500 624.6700 894.5000 627.6700 ;
      RECT 881.2000 624.6700 886.3500 627.6700 ;
      RECT 873.0500 624.6700 878.2000 627.6700 ;
      RECT 864.9000 624.6700 870.0500 627.6700 ;
      RECT 856.7500 624.6700 861.9000 627.6700 ;
      RECT 848.6000 624.6700 853.7500 627.6700 ;
      RECT 840.4500 624.6700 845.6000 627.6700 ;
      RECT 832.3000 624.6700 837.4500 627.6700 ;
      RECT 824.1500 624.6700 829.3000 627.6700 ;
      RECT 816.0000 624.6700 821.1500 627.6700 ;
      RECT 807.8500 624.6700 813.0000 627.6700 ;
      RECT 799.7000 624.6700 804.8500 627.6700 ;
      RECT 791.5500 624.6700 796.7000 627.6700 ;
      RECT 783.4000 624.6700 788.5500 627.6700 ;
      RECT 775.2500 624.6700 780.4000 627.6700 ;
      RECT 767.1000 624.6700 772.2500 627.6700 ;
      RECT 758.9500 624.6700 764.1000 627.6700 ;
      RECT 750.8000 624.6700 755.9500 627.6700 ;
      RECT 742.6500 624.6700 747.8000 627.6700 ;
      RECT 734.5000 624.6700 739.6500 627.6700 ;
      RECT 726.3500 624.6700 731.5000 627.6700 ;
      RECT 718.2000 624.6700 723.3500 627.6700 ;
      RECT 710.0500 624.6700 715.2000 627.6700 ;
      RECT 701.9000 624.6700 707.0500 627.6700 ;
      RECT 693.7500 624.6700 698.9000 627.6700 ;
      RECT 685.6000 624.6700 690.7500 627.6700 ;
      RECT 677.4500 624.6700 682.6000 627.6700 ;
      RECT 669.3000 624.6700 674.4500 627.6700 ;
      RECT 661.1500 624.6700 666.3000 627.6700 ;
      RECT 653.0000 624.6700 658.1500 627.6700 ;
      RECT 644.8500 624.6700 650.0000 627.6700 ;
      RECT 636.7000 624.6700 641.8500 627.6700 ;
      RECT 628.5500 624.6700 633.7000 627.6700 ;
      RECT 620.4000 624.6700 625.5500 627.6700 ;
      RECT 612.2500 624.6700 617.4000 627.6700 ;
      RECT 604.1000 624.6700 609.2500 627.6700 ;
      RECT 595.9500 624.6700 601.1000 627.6700 ;
      RECT 587.8000 624.6700 592.9500 627.6700 ;
      RECT 579.6500 624.6700 584.8000 627.6700 ;
      RECT 571.5000 624.6700 576.6500 627.6700 ;
      RECT 563.3500 624.6700 568.5000 627.6700 ;
      RECT 555.2000 624.6700 560.3500 627.6700 ;
      RECT 547.0500 624.6700 552.2000 627.6700 ;
      RECT 538.9000 624.6700 544.0500 627.6700 ;
      RECT 530.7500 624.6700 535.9000 627.6700 ;
      RECT 522.6000 624.6700 527.7500 627.6700 ;
      RECT 514.4500 624.6700 519.6000 627.6700 ;
      RECT 506.3000 624.6700 511.4500 627.6700 ;
      RECT 498.1500 624.6700 503.3000 627.6700 ;
      RECT 490.0000 624.6700 495.1500 627.6700 ;
      RECT 481.8500 624.6700 487.0000 627.6700 ;
      RECT 473.7000 624.6700 478.8500 627.6700 ;
      RECT 465.5500 624.6700 470.7000 627.6700 ;
      RECT 457.4000 624.6700 462.5500 627.6700 ;
      RECT 449.2500 624.6700 454.4000 627.6700 ;
      RECT 441.1000 624.6700 446.2500 627.6700 ;
      RECT 432.9500 624.6700 438.1000 627.6700 ;
      RECT 424.8000 624.6700 429.9500 627.6700 ;
      RECT 416.6500 624.6700 421.8000 627.6700 ;
      RECT 396.5000 624.6700 413.6500 627.6700 ;
      RECT 346.5000 624.6700 393.5000 627.6700 ;
      RECT 326.4650 624.6700 343.5000 627.6700 ;
      RECT 317.9500 624.6700 323.4650 627.6700 ;
      RECT 309.4350 624.6700 314.9500 627.6700 ;
      RECT 300.9200 624.6700 306.4350 627.6700 ;
      RECT 292.4050 624.6700 297.9200 627.6700 ;
      RECT 283.8900 624.6700 289.4050 627.6700 ;
      RECT 275.3750 624.6700 280.8900 627.6700 ;
      RECT 266.8600 624.6700 272.3750 627.6700 ;
      RECT 258.3450 624.6700 263.8600 627.6700 ;
      RECT 249.8300 624.6700 255.3450 627.6700 ;
      RECT 241.3150 624.6700 246.8300 627.6700 ;
      RECT 232.8000 624.6700 238.3150 627.6700 ;
      RECT 224.2850 624.6700 229.8000 627.6700 ;
      RECT 215.7700 624.6700 221.2850 627.6700 ;
      RECT 207.2550 624.6700 212.7700 627.6700 ;
      RECT 198.7400 624.6700 204.2550 627.6700 ;
      RECT 190.2250 624.6700 195.7400 627.6700 ;
      RECT 181.7100 624.6700 187.2250 627.6700 ;
      RECT 173.1950 624.6700 178.7100 627.6700 ;
      RECT 164.6800 624.6700 170.1950 627.6700 ;
      RECT 156.1650 624.6700 161.6800 627.6700 ;
      RECT 147.6500 624.6700 153.1650 627.6700 ;
      RECT 139.1350 624.6700 144.6500 627.6700 ;
      RECT 130.6200 624.6700 136.1350 627.6700 ;
      RECT 122.1050 624.6700 127.6200 627.6700 ;
      RECT 113.5900 624.6700 119.1050 627.6700 ;
      RECT 105.0750 624.6700 110.5900 627.6700 ;
      RECT 96.5600 624.6700 102.0750 627.6700 ;
      RECT 88.0450 624.6700 93.5600 627.6700 ;
      RECT 79.5300 624.6700 85.0450 627.6700 ;
      RECT 71.0150 624.6700 76.5300 627.6700 ;
      RECT 62.5000 624.6700 68.0150 627.6700 ;
      RECT 46.5000 624.6700 59.5000 627.6700 ;
      RECT 8.5000 624.6700 43.5000 627.6700 ;
      RECT 0.0000 624.6700 5.5000 627.6700 ;
      RECT 0.0000 623.1000 1120.0000 624.6700 ;
      RECT 1116.6000 622.6700 1120.0000 623.1000 ;
      RECT 0.0000 620.5750 1113.6000 623.1000 ;
      RECT 1118.5000 619.6700 1120.0000 622.6700 ;
      RECT 1114.5000 617.5750 1120.0000 619.6700 ;
      RECT 1076.5000 617.5750 1111.5000 620.5750 ;
      RECT 1060.5000 617.5750 1073.5000 620.5750 ;
      RECT 1052.3500 617.5750 1057.5000 620.5750 ;
      RECT 1044.2000 617.5750 1049.3500 620.5750 ;
      RECT 1036.0500 617.5750 1041.2000 620.5750 ;
      RECT 1027.9000 617.5750 1033.0500 620.5750 ;
      RECT 1019.7500 617.5750 1024.9000 620.5750 ;
      RECT 1011.6000 617.5750 1016.7500 620.5750 ;
      RECT 1003.4500 617.5750 1008.6000 620.5750 ;
      RECT 995.3000 617.5750 1000.4500 620.5750 ;
      RECT 987.1500 617.5750 992.3000 620.5750 ;
      RECT 979.0000 617.5750 984.1500 620.5750 ;
      RECT 970.8500 617.5750 976.0000 620.5750 ;
      RECT 962.7000 617.5750 967.8500 620.5750 ;
      RECT 954.5500 617.5750 959.7000 620.5750 ;
      RECT 946.4000 617.5750 951.5500 620.5750 ;
      RECT 938.2500 617.5750 943.4000 620.5750 ;
      RECT 930.1000 617.5750 935.2500 620.5750 ;
      RECT 921.9500 617.5750 927.1000 620.5750 ;
      RECT 913.8000 617.5750 918.9500 620.5750 ;
      RECT 905.6500 617.5750 910.8000 620.5750 ;
      RECT 897.5000 617.5750 902.6500 620.5750 ;
      RECT 889.3500 617.5750 894.5000 620.5750 ;
      RECT 881.2000 617.5750 886.3500 620.5750 ;
      RECT 873.0500 617.5750 878.2000 620.5750 ;
      RECT 864.9000 617.5750 870.0500 620.5750 ;
      RECT 856.7500 617.5750 861.9000 620.5750 ;
      RECT 848.6000 617.5750 853.7500 620.5750 ;
      RECT 840.4500 617.5750 845.6000 620.5750 ;
      RECT 832.3000 617.5750 837.4500 620.5750 ;
      RECT 824.1500 617.5750 829.3000 620.5750 ;
      RECT 816.0000 617.5750 821.1500 620.5750 ;
      RECT 807.8500 617.5750 813.0000 620.5750 ;
      RECT 799.7000 617.5750 804.8500 620.5750 ;
      RECT 791.5500 617.5750 796.7000 620.5750 ;
      RECT 783.4000 617.5750 788.5500 620.5750 ;
      RECT 775.2500 617.5750 780.4000 620.5750 ;
      RECT 767.1000 617.5750 772.2500 620.5750 ;
      RECT 758.9500 617.5750 764.1000 620.5750 ;
      RECT 750.8000 617.5750 755.9500 620.5750 ;
      RECT 742.6500 617.5750 747.8000 620.5750 ;
      RECT 734.5000 617.5750 739.6500 620.5750 ;
      RECT 726.3500 617.5750 731.5000 620.5750 ;
      RECT 718.2000 617.5750 723.3500 620.5750 ;
      RECT 710.0500 617.5750 715.2000 620.5750 ;
      RECT 701.9000 617.5750 707.0500 620.5750 ;
      RECT 693.7500 617.5750 698.9000 620.5750 ;
      RECT 685.6000 617.5750 690.7500 620.5750 ;
      RECT 677.4500 617.5750 682.6000 620.5750 ;
      RECT 669.3000 617.5750 674.4500 620.5750 ;
      RECT 661.1500 617.5750 666.3000 620.5750 ;
      RECT 653.0000 617.5750 658.1500 620.5750 ;
      RECT 644.8500 617.5750 650.0000 620.5750 ;
      RECT 636.7000 617.5750 641.8500 620.5750 ;
      RECT 628.5500 617.5750 633.7000 620.5750 ;
      RECT 620.4000 617.5750 625.5500 620.5750 ;
      RECT 612.2500 617.5750 617.4000 620.5750 ;
      RECT 604.1000 617.5750 609.2500 620.5750 ;
      RECT 595.9500 617.5750 601.1000 620.5750 ;
      RECT 587.8000 617.5750 592.9500 620.5750 ;
      RECT 579.6500 617.5750 584.8000 620.5750 ;
      RECT 571.5000 617.5750 576.6500 620.5750 ;
      RECT 563.3500 617.5750 568.5000 620.5750 ;
      RECT 555.2000 617.5750 560.3500 620.5750 ;
      RECT 547.0500 617.5750 552.2000 620.5750 ;
      RECT 538.9000 617.5750 544.0500 620.5750 ;
      RECT 530.7500 617.5750 535.9000 620.5750 ;
      RECT 522.6000 617.5750 527.7500 620.5750 ;
      RECT 514.4500 617.5750 519.6000 620.5750 ;
      RECT 506.3000 617.5750 511.4500 620.5750 ;
      RECT 498.1500 617.5750 503.3000 620.5750 ;
      RECT 490.0000 617.5750 495.1500 620.5750 ;
      RECT 481.8500 617.5750 487.0000 620.5750 ;
      RECT 473.7000 617.5750 478.8500 620.5750 ;
      RECT 465.5500 617.5750 470.7000 620.5750 ;
      RECT 457.4000 617.5750 462.5500 620.5750 ;
      RECT 449.2500 617.5750 454.4000 620.5750 ;
      RECT 441.1000 617.5750 446.2500 620.5750 ;
      RECT 432.9500 617.5750 438.1000 620.5750 ;
      RECT 424.8000 617.5750 429.9500 620.5750 ;
      RECT 416.6500 617.5750 421.8000 620.5750 ;
      RECT 396.5000 617.5750 413.6500 620.5750 ;
      RECT 346.5000 617.5750 393.5000 620.5750 ;
      RECT 326.4650 617.5750 343.5000 620.5750 ;
      RECT 317.9500 617.5750 323.4650 620.5750 ;
      RECT 309.4350 617.5750 314.9500 620.5750 ;
      RECT 300.9200 617.5750 306.4350 620.5750 ;
      RECT 292.4050 617.5750 297.9200 620.5750 ;
      RECT 283.8900 617.5750 289.4050 620.5750 ;
      RECT 275.3750 617.5750 280.8900 620.5750 ;
      RECT 266.8600 617.5750 272.3750 620.5750 ;
      RECT 258.3450 617.5750 263.8600 620.5750 ;
      RECT 249.8300 617.5750 255.3450 620.5750 ;
      RECT 241.3150 617.5750 246.8300 620.5750 ;
      RECT 232.8000 617.5750 238.3150 620.5750 ;
      RECT 224.2850 617.5750 229.8000 620.5750 ;
      RECT 215.7700 617.5750 221.2850 620.5750 ;
      RECT 207.2550 617.5750 212.7700 620.5750 ;
      RECT 198.7400 617.5750 204.2550 620.5750 ;
      RECT 190.2250 617.5750 195.7400 620.5750 ;
      RECT 181.7100 617.5750 187.2250 620.5750 ;
      RECT 173.1950 617.5750 178.7100 620.5750 ;
      RECT 164.6800 617.5750 170.1950 620.5750 ;
      RECT 156.1650 617.5750 161.6800 620.5750 ;
      RECT 147.6500 617.5750 153.1650 620.5750 ;
      RECT 139.1350 617.5750 144.6500 620.5750 ;
      RECT 130.6200 617.5750 136.1350 620.5750 ;
      RECT 122.1050 617.5750 127.6200 620.5750 ;
      RECT 113.5900 617.5750 119.1050 620.5750 ;
      RECT 105.0750 617.5750 110.5900 620.5750 ;
      RECT 96.5600 617.5750 102.0750 620.5750 ;
      RECT 88.0450 617.5750 93.5600 620.5750 ;
      RECT 79.5300 617.5750 85.0450 620.5750 ;
      RECT 71.0150 617.5750 76.5300 620.5750 ;
      RECT 62.5000 617.5750 68.0150 620.5750 ;
      RECT 46.5000 617.5750 59.5000 620.5750 ;
      RECT 8.5000 617.5750 43.5000 620.5750 ;
      RECT 0.0000 617.5750 5.5000 620.5750 ;
      RECT 0.0000 616.1000 1120.0000 617.5750 ;
      RECT 1116.6000 615.5750 1120.0000 616.1000 ;
      RECT 0.0000 613.4800 1113.6000 616.1000 ;
      RECT 1118.5000 612.5750 1120.0000 615.5750 ;
      RECT 1114.5000 610.4800 1120.0000 612.5750 ;
      RECT 1076.5000 610.4800 1111.5000 613.4800 ;
      RECT 1060.5000 610.4800 1073.5000 613.4800 ;
      RECT 1052.3500 610.4800 1057.5000 613.4800 ;
      RECT 1044.2000 610.4800 1049.3500 613.4800 ;
      RECT 1036.0500 610.4800 1041.2000 613.4800 ;
      RECT 1027.9000 610.4800 1033.0500 613.4800 ;
      RECT 1019.7500 610.4800 1024.9000 613.4800 ;
      RECT 1011.6000 610.4800 1016.7500 613.4800 ;
      RECT 1003.4500 610.4800 1008.6000 613.4800 ;
      RECT 995.3000 610.4800 1000.4500 613.4800 ;
      RECT 987.1500 610.4800 992.3000 613.4800 ;
      RECT 979.0000 610.4800 984.1500 613.4800 ;
      RECT 970.8500 610.4800 976.0000 613.4800 ;
      RECT 962.7000 610.4800 967.8500 613.4800 ;
      RECT 954.5500 610.4800 959.7000 613.4800 ;
      RECT 946.4000 610.4800 951.5500 613.4800 ;
      RECT 938.2500 610.4800 943.4000 613.4800 ;
      RECT 930.1000 610.4800 935.2500 613.4800 ;
      RECT 921.9500 610.4800 927.1000 613.4800 ;
      RECT 913.8000 610.4800 918.9500 613.4800 ;
      RECT 905.6500 610.4800 910.8000 613.4800 ;
      RECT 897.5000 610.4800 902.6500 613.4800 ;
      RECT 889.3500 610.4800 894.5000 613.4800 ;
      RECT 881.2000 610.4800 886.3500 613.4800 ;
      RECT 873.0500 610.4800 878.2000 613.4800 ;
      RECT 864.9000 610.4800 870.0500 613.4800 ;
      RECT 856.7500 610.4800 861.9000 613.4800 ;
      RECT 848.6000 610.4800 853.7500 613.4800 ;
      RECT 840.4500 610.4800 845.6000 613.4800 ;
      RECT 832.3000 610.4800 837.4500 613.4800 ;
      RECT 824.1500 610.4800 829.3000 613.4800 ;
      RECT 816.0000 610.4800 821.1500 613.4800 ;
      RECT 807.8500 610.4800 813.0000 613.4800 ;
      RECT 799.7000 610.4800 804.8500 613.4800 ;
      RECT 791.5500 610.4800 796.7000 613.4800 ;
      RECT 783.4000 610.4800 788.5500 613.4800 ;
      RECT 775.2500 610.4800 780.4000 613.4800 ;
      RECT 767.1000 610.4800 772.2500 613.4800 ;
      RECT 758.9500 610.4800 764.1000 613.4800 ;
      RECT 750.8000 610.4800 755.9500 613.4800 ;
      RECT 742.6500 610.4800 747.8000 613.4800 ;
      RECT 734.5000 610.4800 739.6500 613.4800 ;
      RECT 726.3500 610.4800 731.5000 613.4800 ;
      RECT 718.2000 610.4800 723.3500 613.4800 ;
      RECT 710.0500 610.4800 715.2000 613.4800 ;
      RECT 701.9000 610.4800 707.0500 613.4800 ;
      RECT 693.7500 610.4800 698.9000 613.4800 ;
      RECT 685.6000 610.4800 690.7500 613.4800 ;
      RECT 677.4500 610.4800 682.6000 613.4800 ;
      RECT 669.3000 610.4800 674.4500 613.4800 ;
      RECT 661.1500 610.4800 666.3000 613.4800 ;
      RECT 653.0000 610.4800 658.1500 613.4800 ;
      RECT 644.8500 610.4800 650.0000 613.4800 ;
      RECT 636.7000 610.4800 641.8500 613.4800 ;
      RECT 628.5500 610.4800 633.7000 613.4800 ;
      RECT 620.4000 610.4800 625.5500 613.4800 ;
      RECT 612.2500 610.4800 617.4000 613.4800 ;
      RECT 604.1000 610.4800 609.2500 613.4800 ;
      RECT 595.9500 610.4800 601.1000 613.4800 ;
      RECT 587.8000 610.4800 592.9500 613.4800 ;
      RECT 579.6500 610.4800 584.8000 613.4800 ;
      RECT 571.5000 610.4800 576.6500 613.4800 ;
      RECT 563.3500 610.4800 568.5000 613.4800 ;
      RECT 555.2000 610.4800 560.3500 613.4800 ;
      RECT 547.0500 610.4800 552.2000 613.4800 ;
      RECT 538.9000 610.4800 544.0500 613.4800 ;
      RECT 530.7500 610.4800 535.9000 613.4800 ;
      RECT 522.6000 610.4800 527.7500 613.4800 ;
      RECT 514.4500 610.4800 519.6000 613.4800 ;
      RECT 506.3000 610.4800 511.4500 613.4800 ;
      RECT 498.1500 610.4800 503.3000 613.4800 ;
      RECT 490.0000 610.4800 495.1500 613.4800 ;
      RECT 481.8500 610.4800 487.0000 613.4800 ;
      RECT 473.7000 610.4800 478.8500 613.4800 ;
      RECT 465.5500 610.4800 470.7000 613.4800 ;
      RECT 457.4000 610.4800 462.5500 613.4800 ;
      RECT 449.2500 610.4800 454.4000 613.4800 ;
      RECT 441.1000 610.4800 446.2500 613.4800 ;
      RECT 432.9500 610.4800 438.1000 613.4800 ;
      RECT 424.8000 610.4800 429.9500 613.4800 ;
      RECT 416.6500 610.4800 421.8000 613.4800 ;
      RECT 396.5000 610.4800 413.6500 613.4800 ;
      RECT 346.5000 610.4800 393.5000 613.4800 ;
      RECT 326.4650 610.4800 343.5000 613.4800 ;
      RECT 317.9500 610.4800 323.4650 613.4800 ;
      RECT 309.4350 610.4800 314.9500 613.4800 ;
      RECT 300.9200 610.4800 306.4350 613.4800 ;
      RECT 292.4050 610.4800 297.9200 613.4800 ;
      RECT 283.8900 610.4800 289.4050 613.4800 ;
      RECT 275.3750 610.4800 280.8900 613.4800 ;
      RECT 266.8600 610.4800 272.3750 613.4800 ;
      RECT 258.3450 610.4800 263.8600 613.4800 ;
      RECT 249.8300 610.4800 255.3450 613.4800 ;
      RECT 241.3150 610.4800 246.8300 613.4800 ;
      RECT 232.8000 610.4800 238.3150 613.4800 ;
      RECT 224.2850 610.4800 229.8000 613.4800 ;
      RECT 215.7700 610.4800 221.2850 613.4800 ;
      RECT 207.2550 610.4800 212.7700 613.4800 ;
      RECT 198.7400 610.4800 204.2550 613.4800 ;
      RECT 190.2250 610.4800 195.7400 613.4800 ;
      RECT 181.7100 610.4800 187.2250 613.4800 ;
      RECT 173.1950 610.4800 178.7100 613.4800 ;
      RECT 164.6800 610.4800 170.1950 613.4800 ;
      RECT 156.1650 610.4800 161.6800 613.4800 ;
      RECT 147.6500 610.4800 153.1650 613.4800 ;
      RECT 139.1350 610.4800 144.6500 613.4800 ;
      RECT 130.6200 610.4800 136.1350 613.4800 ;
      RECT 122.1050 610.4800 127.6200 613.4800 ;
      RECT 113.5900 610.4800 119.1050 613.4800 ;
      RECT 105.0750 610.4800 110.5900 613.4800 ;
      RECT 96.5600 610.4800 102.0750 613.4800 ;
      RECT 88.0450 610.4800 93.5600 613.4800 ;
      RECT 79.5300 610.4800 85.0450 613.4800 ;
      RECT 71.0150 610.4800 76.5300 613.4800 ;
      RECT 62.5000 610.4800 68.0150 613.4800 ;
      RECT 46.5000 610.4800 59.5000 613.4800 ;
      RECT 8.5000 610.4800 43.5000 613.4800 ;
      RECT 0.0000 610.4800 5.5000 613.4800 ;
      RECT 0.0000 608.9000 1120.0000 610.4800 ;
      RECT 1116.6000 608.4800 1120.0000 608.9000 ;
      RECT 0.0000 606.3850 1113.6000 608.9000 ;
      RECT 1118.5000 605.4800 1120.0000 608.4800 ;
      RECT 1114.5000 603.3850 1120.0000 605.4800 ;
      RECT 1076.5000 603.3850 1111.5000 606.3850 ;
      RECT 1060.5000 603.3850 1073.5000 606.3850 ;
      RECT 1052.3500 603.3850 1057.5000 606.3850 ;
      RECT 1044.2000 603.3850 1049.3500 606.3850 ;
      RECT 1036.0500 603.3850 1041.2000 606.3850 ;
      RECT 1027.9000 603.3850 1033.0500 606.3850 ;
      RECT 1019.7500 603.3850 1024.9000 606.3850 ;
      RECT 1011.6000 603.3850 1016.7500 606.3850 ;
      RECT 1003.4500 603.3850 1008.6000 606.3850 ;
      RECT 995.3000 603.3850 1000.4500 606.3850 ;
      RECT 987.1500 603.3850 992.3000 606.3850 ;
      RECT 979.0000 603.3850 984.1500 606.3850 ;
      RECT 970.8500 603.3850 976.0000 606.3850 ;
      RECT 962.7000 603.3850 967.8500 606.3850 ;
      RECT 954.5500 603.3850 959.7000 606.3850 ;
      RECT 946.4000 603.3850 951.5500 606.3850 ;
      RECT 938.2500 603.3850 943.4000 606.3850 ;
      RECT 930.1000 603.3850 935.2500 606.3850 ;
      RECT 921.9500 603.3850 927.1000 606.3850 ;
      RECT 913.8000 603.3850 918.9500 606.3850 ;
      RECT 905.6500 603.3850 910.8000 606.3850 ;
      RECT 897.5000 603.3850 902.6500 606.3850 ;
      RECT 889.3500 603.3850 894.5000 606.3850 ;
      RECT 881.2000 603.3850 886.3500 606.3850 ;
      RECT 873.0500 603.3850 878.2000 606.3850 ;
      RECT 864.9000 603.3850 870.0500 606.3850 ;
      RECT 856.7500 603.3850 861.9000 606.3850 ;
      RECT 848.6000 603.3850 853.7500 606.3850 ;
      RECT 840.4500 603.3850 845.6000 606.3850 ;
      RECT 832.3000 603.3850 837.4500 606.3850 ;
      RECT 824.1500 603.3850 829.3000 606.3850 ;
      RECT 816.0000 603.3850 821.1500 606.3850 ;
      RECT 807.8500 603.3850 813.0000 606.3850 ;
      RECT 799.7000 603.3850 804.8500 606.3850 ;
      RECT 791.5500 603.3850 796.7000 606.3850 ;
      RECT 783.4000 603.3850 788.5500 606.3850 ;
      RECT 775.2500 603.3850 780.4000 606.3850 ;
      RECT 767.1000 603.3850 772.2500 606.3850 ;
      RECT 758.9500 603.3850 764.1000 606.3850 ;
      RECT 750.8000 603.3850 755.9500 606.3850 ;
      RECT 742.6500 603.3850 747.8000 606.3850 ;
      RECT 734.5000 603.3850 739.6500 606.3850 ;
      RECT 726.3500 603.3850 731.5000 606.3850 ;
      RECT 718.2000 603.3850 723.3500 606.3850 ;
      RECT 710.0500 603.3850 715.2000 606.3850 ;
      RECT 701.9000 603.3850 707.0500 606.3850 ;
      RECT 693.7500 603.3850 698.9000 606.3850 ;
      RECT 685.6000 603.3850 690.7500 606.3850 ;
      RECT 677.4500 603.3850 682.6000 606.3850 ;
      RECT 669.3000 603.3850 674.4500 606.3850 ;
      RECT 661.1500 603.3850 666.3000 606.3850 ;
      RECT 653.0000 603.3850 658.1500 606.3850 ;
      RECT 644.8500 603.3850 650.0000 606.3850 ;
      RECT 636.7000 603.3850 641.8500 606.3850 ;
      RECT 628.5500 603.3850 633.7000 606.3850 ;
      RECT 620.4000 603.3850 625.5500 606.3850 ;
      RECT 612.2500 603.3850 617.4000 606.3850 ;
      RECT 604.1000 603.3850 609.2500 606.3850 ;
      RECT 595.9500 603.3850 601.1000 606.3850 ;
      RECT 587.8000 603.3850 592.9500 606.3850 ;
      RECT 579.6500 603.3850 584.8000 606.3850 ;
      RECT 571.5000 603.3850 576.6500 606.3850 ;
      RECT 563.3500 603.3850 568.5000 606.3850 ;
      RECT 555.2000 603.3850 560.3500 606.3850 ;
      RECT 547.0500 603.3850 552.2000 606.3850 ;
      RECT 538.9000 603.3850 544.0500 606.3850 ;
      RECT 530.7500 603.3850 535.9000 606.3850 ;
      RECT 522.6000 603.3850 527.7500 606.3850 ;
      RECT 514.4500 603.3850 519.6000 606.3850 ;
      RECT 506.3000 603.3850 511.4500 606.3850 ;
      RECT 498.1500 603.3850 503.3000 606.3850 ;
      RECT 490.0000 603.3850 495.1500 606.3850 ;
      RECT 481.8500 603.3850 487.0000 606.3850 ;
      RECT 473.7000 603.3850 478.8500 606.3850 ;
      RECT 465.5500 603.3850 470.7000 606.3850 ;
      RECT 457.4000 603.3850 462.5500 606.3850 ;
      RECT 449.2500 603.3850 454.4000 606.3850 ;
      RECT 441.1000 603.3850 446.2500 606.3850 ;
      RECT 432.9500 603.3850 438.1000 606.3850 ;
      RECT 424.8000 603.3850 429.9500 606.3850 ;
      RECT 416.6500 603.3850 421.8000 606.3850 ;
      RECT 396.5000 603.3850 413.6500 606.3850 ;
      RECT 346.5000 603.3850 393.5000 606.3850 ;
      RECT 326.4650 603.3850 343.5000 606.3850 ;
      RECT 317.9500 603.3850 323.4650 606.3850 ;
      RECT 309.4350 603.3850 314.9500 606.3850 ;
      RECT 300.9200 603.3850 306.4350 606.3850 ;
      RECT 292.4050 603.3850 297.9200 606.3850 ;
      RECT 283.8900 603.3850 289.4050 606.3850 ;
      RECT 275.3750 603.3850 280.8900 606.3850 ;
      RECT 266.8600 603.3850 272.3750 606.3850 ;
      RECT 258.3450 603.3850 263.8600 606.3850 ;
      RECT 249.8300 603.3850 255.3450 606.3850 ;
      RECT 241.3150 603.3850 246.8300 606.3850 ;
      RECT 232.8000 603.3850 238.3150 606.3850 ;
      RECT 224.2850 603.3850 229.8000 606.3850 ;
      RECT 215.7700 603.3850 221.2850 606.3850 ;
      RECT 207.2550 603.3850 212.7700 606.3850 ;
      RECT 198.7400 603.3850 204.2550 606.3850 ;
      RECT 190.2250 603.3850 195.7400 606.3850 ;
      RECT 181.7100 603.3850 187.2250 606.3850 ;
      RECT 173.1950 603.3850 178.7100 606.3850 ;
      RECT 164.6800 603.3850 170.1950 606.3850 ;
      RECT 156.1650 603.3850 161.6800 606.3850 ;
      RECT 147.6500 603.3850 153.1650 606.3850 ;
      RECT 139.1350 603.3850 144.6500 606.3850 ;
      RECT 130.6200 603.3850 136.1350 606.3850 ;
      RECT 122.1050 603.3850 127.6200 606.3850 ;
      RECT 113.5900 603.3850 119.1050 606.3850 ;
      RECT 105.0750 603.3850 110.5900 606.3850 ;
      RECT 96.5600 603.3850 102.0750 606.3850 ;
      RECT 88.0450 603.3850 93.5600 606.3850 ;
      RECT 79.5300 603.3850 85.0450 606.3850 ;
      RECT 71.0150 603.3850 76.5300 606.3850 ;
      RECT 62.5000 603.3850 68.0150 606.3850 ;
      RECT 46.5000 603.3850 59.5000 606.3850 ;
      RECT 8.5000 603.3850 43.5000 606.3850 ;
      RECT 0.0000 603.3850 5.5000 606.3850 ;
      RECT 0.0000 601.9000 1120.0000 603.3850 ;
      RECT 1116.6000 601.3850 1120.0000 601.9000 ;
      RECT 0.0000 599.2900 1113.6000 601.9000 ;
      RECT 1118.5000 598.3850 1120.0000 601.3850 ;
      RECT 1114.5000 596.2900 1120.0000 598.3850 ;
      RECT 1076.5000 596.2900 1111.5000 599.2900 ;
      RECT 1060.5000 596.2900 1073.5000 599.2900 ;
      RECT 1052.3500 596.2900 1057.5000 599.2900 ;
      RECT 1044.2000 596.2900 1049.3500 599.2900 ;
      RECT 1036.0500 596.2900 1041.2000 599.2900 ;
      RECT 1027.9000 596.2900 1033.0500 599.2900 ;
      RECT 1019.7500 596.2900 1024.9000 599.2900 ;
      RECT 1011.6000 596.2900 1016.7500 599.2900 ;
      RECT 1003.4500 596.2900 1008.6000 599.2900 ;
      RECT 995.3000 596.2900 1000.4500 599.2900 ;
      RECT 987.1500 596.2900 992.3000 599.2900 ;
      RECT 979.0000 596.2900 984.1500 599.2900 ;
      RECT 970.8500 596.2900 976.0000 599.2900 ;
      RECT 962.7000 596.2900 967.8500 599.2900 ;
      RECT 954.5500 596.2900 959.7000 599.2900 ;
      RECT 946.4000 596.2900 951.5500 599.2900 ;
      RECT 938.2500 596.2900 943.4000 599.2900 ;
      RECT 930.1000 596.2900 935.2500 599.2900 ;
      RECT 921.9500 596.2900 927.1000 599.2900 ;
      RECT 913.8000 596.2900 918.9500 599.2900 ;
      RECT 905.6500 596.2900 910.8000 599.2900 ;
      RECT 897.5000 596.2900 902.6500 599.2900 ;
      RECT 889.3500 596.2900 894.5000 599.2900 ;
      RECT 881.2000 596.2900 886.3500 599.2900 ;
      RECT 873.0500 596.2900 878.2000 599.2900 ;
      RECT 864.9000 596.2900 870.0500 599.2900 ;
      RECT 856.7500 596.2900 861.9000 599.2900 ;
      RECT 848.6000 596.2900 853.7500 599.2900 ;
      RECT 840.4500 596.2900 845.6000 599.2900 ;
      RECT 832.3000 596.2900 837.4500 599.2900 ;
      RECT 824.1500 596.2900 829.3000 599.2900 ;
      RECT 816.0000 596.2900 821.1500 599.2900 ;
      RECT 807.8500 596.2900 813.0000 599.2900 ;
      RECT 799.7000 596.2900 804.8500 599.2900 ;
      RECT 791.5500 596.2900 796.7000 599.2900 ;
      RECT 783.4000 596.2900 788.5500 599.2900 ;
      RECT 775.2500 596.2900 780.4000 599.2900 ;
      RECT 767.1000 596.2900 772.2500 599.2900 ;
      RECT 758.9500 596.2900 764.1000 599.2900 ;
      RECT 750.8000 596.2900 755.9500 599.2900 ;
      RECT 742.6500 596.2900 747.8000 599.2900 ;
      RECT 734.5000 596.2900 739.6500 599.2900 ;
      RECT 726.3500 596.2900 731.5000 599.2900 ;
      RECT 718.2000 596.2900 723.3500 599.2900 ;
      RECT 710.0500 596.2900 715.2000 599.2900 ;
      RECT 701.9000 596.2900 707.0500 599.2900 ;
      RECT 693.7500 596.2900 698.9000 599.2900 ;
      RECT 685.6000 596.2900 690.7500 599.2900 ;
      RECT 677.4500 596.2900 682.6000 599.2900 ;
      RECT 669.3000 596.2900 674.4500 599.2900 ;
      RECT 661.1500 596.2900 666.3000 599.2900 ;
      RECT 653.0000 596.2900 658.1500 599.2900 ;
      RECT 644.8500 596.2900 650.0000 599.2900 ;
      RECT 636.7000 596.2900 641.8500 599.2900 ;
      RECT 628.5500 596.2900 633.7000 599.2900 ;
      RECT 620.4000 596.2900 625.5500 599.2900 ;
      RECT 612.2500 596.2900 617.4000 599.2900 ;
      RECT 604.1000 596.2900 609.2500 599.2900 ;
      RECT 595.9500 596.2900 601.1000 599.2900 ;
      RECT 587.8000 596.2900 592.9500 599.2900 ;
      RECT 579.6500 596.2900 584.8000 599.2900 ;
      RECT 571.5000 596.2900 576.6500 599.2900 ;
      RECT 563.3500 596.2900 568.5000 599.2900 ;
      RECT 555.2000 596.2900 560.3500 599.2900 ;
      RECT 547.0500 596.2900 552.2000 599.2900 ;
      RECT 538.9000 596.2900 544.0500 599.2900 ;
      RECT 530.7500 596.2900 535.9000 599.2900 ;
      RECT 522.6000 596.2900 527.7500 599.2900 ;
      RECT 514.4500 596.2900 519.6000 599.2900 ;
      RECT 506.3000 596.2900 511.4500 599.2900 ;
      RECT 498.1500 596.2900 503.3000 599.2900 ;
      RECT 490.0000 596.2900 495.1500 599.2900 ;
      RECT 481.8500 596.2900 487.0000 599.2900 ;
      RECT 473.7000 596.2900 478.8500 599.2900 ;
      RECT 465.5500 596.2900 470.7000 599.2900 ;
      RECT 457.4000 596.2900 462.5500 599.2900 ;
      RECT 449.2500 596.2900 454.4000 599.2900 ;
      RECT 441.1000 596.2900 446.2500 599.2900 ;
      RECT 432.9500 596.2900 438.1000 599.2900 ;
      RECT 424.8000 596.2900 429.9500 599.2900 ;
      RECT 416.6500 596.2900 421.8000 599.2900 ;
      RECT 396.5000 596.2900 413.6500 599.2900 ;
      RECT 346.5000 596.2900 393.5000 599.2900 ;
      RECT 326.4650 596.2900 343.5000 599.2900 ;
      RECT 317.9500 596.2900 323.4650 599.2900 ;
      RECT 309.4350 596.2900 314.9500 599.2900 ;
      RECT 300.9200 596.2900 306.4350 599.2900 ;
      RECT 292.4050 596.2900 297.9200 599.2900 ;
      RECT 283.8900 596.2900 289.4050 599.2900 ;
      RECT 275.3750 596.2900 280.8900 599.2900 ;
      RECT 266.8600 596.2900 272.3750 599.2900 ;
      RECT 258.3450 596.2900 263.8600 599.2900 ;
      RECT 249.8300 596.2900 255.3450 599.2900 ;
      RECT 241.3150 596.2900 246.8300 599.2900 ;
      RECT 232.8000 596.2900 238.3150 599.2900 ;
      RECT 224.2850 596.2900 229.8000 599.2900 ;
      RECT 215.7700 596.2900 221.2850 599.2900 ;
      RECT 207.2550 596.2900 212.7700 599.2900 ;
      RECT 198.7400 596.2900 204.2550 599.2900 ;
      RECT 190.2250 596.2900 195.7400 599.2900 ;
      RECT 181.7100 596.2900 187.2250 599.2900 ;
      RECT 173.1950 596.2900 178.7100 599.2900 ;
      RECT 164.6800 596.2900 170.1950 599.2900 ;
      RECT 156.1650 596.2900 161.6800 599.2900 ;
      RECT 147.6500 596.2900 153.1650 599.2900 ;
      RECT 139.1350 596.2900 144.6500 599.2900 ;
      RECT 130.6200 596.2900 136.1350 599.2900 ;
      RECT 122.1050 596.2900 127.6200 599.2900 ;
      RECT 113.5900 596.2900 119.1050 599.2900 ;
      RECT 105.0750 596.2900 110.5900 599.2900 ;
      RECT 96.5600 596.2900 102.0750 599.2900 ;
      RECT 88.0450 596.2900 93.5600 599.2900 ;
      RECT 79.5300 596.2900 85.0450 599.2900 ;
      RECT 71.0150 596.2900 76.5300 599.2900 ;
      RECT 62.5000 596.2900 68.0150 599.2900 ;
      RECT 46.5000 596.2900 59.5000 599.2900 ;
      RECT 8.5000 596.2900 43.5000 599.2900 ;
      RECT 0.0000 596.2900 5.5000 599.2900 ;
      RECT 0.0000 594.7000 1120.0000 596.2900 ;
      RECT 1116.6000 594.2900 1120.0000 594.7000 ;
      RECT 0.0000 592.1950 1113.6000 594.7000 ;
      RECT 1118.5000 591.2900 1120.0000 594.2900 ;
      RECT 1114.5000 589.1950 1120.0000 591.2900 ;
      RECT 1076.5000 589.1950 1111.5000 592.1950 ;
      RECT 1060.5000 589.1950 1073.5000 592.1950 ;
      RECT 1052.3500 589.1950 1057.5000 592.1950 ;
      RECT 1044.2000 589.1950 1049.3500 592.1950 ;
      RECT 1036.0500 589.1950 1041.2000 592.1950 ;
      RECT 1027.9000 589.1950 1033.0500 592.1950 ;
      RECT 1019.7500 589.1950 1024.9000 592.1950 ;
      RECT 1011.6000 589.1950 1016.7500 592.1950 ;
      RECT 1003.4500 589.1950 1008.6000 592.1950 ;
      RECT 995.3000 589.1950 1000.4500 592.1950 ;
      RECT 987.1500 589.1950 992.3000 592.1950 ;
      RECT 979.0000 589.1950 984.1500 592.1950 ;
      RECT 970.8500 589.1950 976.0000 592.1950 ;
      RECT 962.7000 589.1950 967.8500 592.1950 ;
      RECT 954.5500 589.1950 959.7000 592.1950 ;
      RECT 946.4000 589.1950 951.5500 592.1950 ;
      RECT 938.2500 589.1950 943.4000 592.1950 ;
      RECT 930.1000 589.1950 935.2500 592.1950 ;
      RECT 921.9500 589.1950 927.1000 592.1950 ;
      RECT 913.8000 589.1950 918.9500 592.1950 ;
      RECT 905.6500 589.1950 910.8000 592.1950 ;
      RECT 897.5000 589.1950 902.6500 592.1950 ;
      RECT 889.3500 589.1950 894.5000 592.1950 ;
      RECT 881.2000 589.1950 886.3500 592.1950 ;
      RECT 873.0500 589.1950 878.2000 592.1950 ;
      RECT 864.9000 589.1950 870.0500 592.1950 ;
      RECT 856.7500 589.1950 861.9000 592.1950 ;
      RECT 848.6000 589.1950 853.7500 592.1950 ;
      RECT 840.4500 589.1950 845.6000 592.1950 ;
      RECT 832.3000 589.1950 837.4500 592.1950 ;
      RECT 824.1500 589.1950 829.3000 592.1950 ;
      RECT 816.0000 589.1950 821.1500 592.1950 ;
      RECT 807.8500 589.1950 813.0000 592.1950 ;
      RECT 799.7000 589.1950 804.8500 592.1950 ;
      RECT 791.5500 589.1950 796.7000 592.1950 ;
      RECT 783.4000 589.1950 788.5500 592.1950 ;
      RECT 775.2500 589.1950 780.4000 592.1950 ;
      RECT 767.1000 589.1950 772.2500 592.1950 ;
      RECT 758.9500 589.1950 764.1000 592.1950 ;
      RECT 750.8000 589.1950 755.9500 592.1950 ;
      RECT 742.6500 589.1950 747.8000 592.1950 ;
      RECT 734.5000 589.1950 739.6500 592.1950 ;
      RECT 726.3500 589.1950 731.5000 592.1950 ;
      RECT 718.2000 589.1950 723.3500 592.1950 ;
      RECT 710.0500 589.1950 715.2000 592.1950 ;
      RECT 701.9000 589.1950 707.0500 592.1950 ;
      RECT 693.7500 589.1950 698.9000 592.1950 ;
      RECT 685.6000 589.1950 690.7500 592.1950 ;
      RECT 677.4500 589.1950 682.6000 592.1950 ;
      RECT 669.3000 589.1950 674.4500 592.1950 ;
      RECT 661.1500 589.1950 666.3000 592.1950 ;
      RECT 653.0000 589.1950 658.1500 592.1950 ;
      RECT 644.8500 589.1950 650.0000 592.1950 ;
      RECT 636.7000 589.1950 641.8500 592.1950 ;
      RECT 628.5500 589.1950 633.7000 592.1950 ;
      RECT 620.4000 589.1950 625.5500 592.1950 ;
      RECT 612.2500 589.1950 617.4000 592.1950 ;
      RECT 604.1000 589.1950 609.2500 592.1950 ;
      RECT 595.9500 589.1950 601.1000 592.1950 ;
      RECT 587.8000 589.1950 592.9500 592.1950 ;
      RECT 579.6500 589.1950 584.8000 592.1950 ;
      RECT 571.5000 589.1950 576.6500 592.1950 ;
      RECT 563.3500 589.1950 568.5000 592.1950 ;
      RECT 555.2000 589.1950 560.3500 592.1950 ;
      RECT 547.0500 589.1950 552.2000 592.1950 ;
      RECT 538.9000 589.1950 544.0500 592.1950 ;
      RECT 530.7500 589.1950 535.9000 592.1950 ;
      RECT 522.6000 589.1950 527.7500 592.1950 ;
      RECT 514.4500 589.1950 519.6000 592.1950 ;
      RECT 506.3000 589.1950 511.4500 592.1950 ;
      RECT 498.1500 589.1950 503.3000 592.1950 ;
      RECT 490.0000 589.1950 495.1500 592.1950 ;
      RECT 481.8500 589.1950 487.0000 592.1950 ;
      RECT 473.7000 589.1950 478.8500 592.1950 ;
      RECT 465.5500 589.1950 470.7000 592.1950 ;
      RECT 457.4000 589.1950 462.5500 592.1950 ;
      RECT 449.2500 589.1950 454.4000 592.1950 ;
      RECT 441.1000 589.1950 446.2500 592.1950 ;
      RECT 432.9500 589.1950 438.1000 592.1950 ;
      RECT 424.8000 589.1950 429.9500 592.1950 ;
      RECT 416.6500 589.1950 421.8000 592.1950 ;
      RECT 396.5000 589.1950 413.6500 592.1950 ;
      RECT 346.5000 589.1950 393.5000 592.1950 ;
      RECT 326.4650 589.1950 343.5000 592.1950 ;
      RECT 317.9500 589.1950 323.4650 592.1950 ;
      RECT 309.4350 589.1950 314.9500 592.1950 ;
      RECT 300.9200 589.1950 306.4350 592.1950 ;
      RECT 292.4050 589.1950 297.9200 592.1950 ;
      RECT 283.8900 589.1950 289.4050 592.1950 ;
      RECT 275.3750 589.1950 280.8900 592.1950 ;
      RECT 266.8600 589.1950 272.3750 592.1950 ;
      RECT 258.3450 589.1950 263.8600 592.1950 ;
      RECT 249.8300 589.1950 255.3450 592.1950 ;
      RECT 241.3150 589.1950 246.8300 592.1950 ;
      RECT 232.8000 589.1950 238.3150 592.1950 ;
      RECT 224.2850 589.1950 229.8000 592.1950 ;
      RECT 215.7700 589.1950 221.2850 592.1950 ;
      RECT 207.2550 589.1950 212.7700 592.1950 ;
      RECT 198.7400 589.1950 204.2550 592.1950 ;
      RECT 190.2250 589.1950 195.7400 592.1950 ;
      RECT 181.7100 589.1950 187.2250 592.1950 ;
      RECT 173.1950 589.1950 178.7100 592.1950 ;
      RECT 164.6800 589.1950 170.1950 592.1950 ;
      RECT 156.1650 589.1950 161.6800 592.1950 ;
      RECT 147.6500 589.1950 153.1650 592.1950 ;
      RECT 139.1350 589.1950 144.6500 592.1950 ;
      RECT 130.6200 589.1950 136.1350 592.1950 ;
      RECT 122.1050 589.1950 127.6200 592.1950 ;
      RECT 113.5900 589.1950 119.1050 592.1950 ;
      RECT 105.0750 589.1950 110.5900 592.1950 ;
      RECT 96.5600 589.1950 102.0750 592.1950 ;
      RECT 88.0450 589.1950 93.5600 592.1950 ;
      RECT 79.5300 589.1950 85.0450 592.1950 ;
      RECT 71.0150 589.1950 76.5300 592.1950 ;
      RECT 62.5000 589.1950 68.0150 592.1950 ;
      RECT 46.5000 589.1950 59.5000 592.1950 ;
      RECT 8.5000 589.1950 43.5000 592.1950 ;
      RECT 0.0000 589.1950 5.5000 592.1950 ;
      RECT 0.0000 587.7000 1120.0000 589.1950 ;
      RECT 1116.6000 587.1950 1120.0000 587.7000 ;
      RECT 0.0000 585.1000 1113.6000 587.7000 ;
      RECT 1118.5000 584.1950 1120.0000 587.1950 ;
      RECT 1114.5000 582.1000 1120.0000 584.1950 ;
      RECT 1076.5000 582.1000 1111.5000 585.1000 ;
      RECT 1060.5000 582.1000 1073.5000 585.1000 ;
      RECT 1052.3500 582.1000 1057.5000 585.1000 ;
      RECT 1044.2000 582.1000 1049.3500 585.1000 ;
      RECT 1036.0500 582.1000 1041.2000 585.1000 ;
      RECT 1027.9000 582.1000 1033.0500 585.1000 ;
      RECT 1019.7500 582.1000 1024.9000 585.1000 ;
      RECT 1011.6000 582.1000 1016.7500 585.1000 ;
      RECT 1003.4500 582.1000 1008.6000 585.1000 ;
      RECT 995.3000 582.1000 1000.4500 585.1000 ;
      RECT 987.1500 582.1000 992.3000 585.1000 ;
      RECT 979.0000 582.1000 984.1500 585.1000 ;
      RECT 970.8500 582.1000 976.0000 585.1000 ;
      RECT 962.7000 582.1000 967.8500 585.1000 ;
      RECT 954.5500 582.1000 959.7000 585.1000 ;
      RECT 946.4000 582.1000 951.5500 585.1000 ;
      RECT 938.2500 582.1000 943.4000 585.1000 ;
      RECT 930.1000 582.1000 935.2500 585.1000 ;
      RECT 921.9500 582.1000 927.1000 585.1000 ;
      RECT 913.8000 582.1000 918.9500 585.1000 ;
      RECT 905.6500 582.1000 910.8000 585.1000 ;
      RECT 897.5000 582.1000 902.6500 585.1000 ;
      RECT 889.3500 582.1000 894.5000 585.1000 ;
      RECT 881.2000 582.1000 886.3500 585.1000 ;
      RECT 873.0500 582.1000 878.2000 585.1000 ;
      RECT 864.9000 582.1000 870.0500 585.1000 ;
      RECT 856.7500 582.1000 861.9000 585.1000 ;
      RECT 848.6000 582.1000 853.7500 585.1000 ;
      RECT 840.4500 582.1000 845.6000 585.1000 ;
      RECT 832.3000 582.1000 837.4500 585.1000 ;
      RECT 824.1500 582.1000 829.3000 585.1000 ;
      RECT 816.0000 582.1000 821.1500 585.1000 ;
      RECT 807.8500 582.1000 813.0000 585.1000 ;
      RECT 799.7000 582.1000 804.8500 585.1000 ;
      RECT 791.5500 582.1000 796.7000 585.1000 ;
      RECT 783.4000 582.1000 788.5500 585.1000 ;
      RECT 775.2500 582.1000 780.4000 585.1000 ;
      RECT 767.1000 582.1000 772.2500 585.1000 ;
      RECT 758.9500 582.1000 764.1000 585.1000 ;
      RECT 750.8000 582.1000 755.9500 585.1000 ;
      RECT 742.6500 582.1000 747.8000 585.1000 ;
      RECT 734.5000 582.1000 739.6500 585.1000 ;
      RECT 726.3500 582.1000 731.5000 585.1000 ;
      RECT 718.2000 582.1000 723.3500 585.1000 ;
      RECT 710.0500 582.1000 715.2000 585.1000 ;
      RECT 701.9000 582.1000 707.0500 585.1000 ;
      RECT 693.7500 582.1000 698.9000 585.1000 ;
      RECT 685.6000 582.1000 690.7500 585.1000 ;
      RECT 677.4500 582.1000 682.6000 585.1000 ;
      RECT 669.3000 582.1000 674.4500 585.1000 ;
      RECT 661.1500 582.1000 666.3000 585.1000 ;
      RECT 653.0000 582.1000 658.1500 585.1000 ;
      RECT 644.8500 582.1000 650.0000 585.1000 ;
      RECT 636.7000 582.1000 641.8500 585.1000 ;
      RECT 628.5500 582.1000 633.7000 585.1000 ;
      RECT 620.4000 582.1000 625.5500 585.1000 ;
      RECT 612.2500 582.1000 617.4000 585.1000 ;
      RECT 604.1000 582.1000 609.2500 585.1000 ;
      RECT 595.9500 582.1000 601.1000 585.1000 ;
      RECT 587.8000 582.1000 592.9500 585.1000 ;
      RECT 579.6500 582.1000 584.8000 585.1000 ;
      RECT 571.5000 582.1000 576.6500 585.1000 ;
      RECT 563.3500 582.1000 568.5000 585.1000 ;
      RECT 555.2000 582.1000 560.3500 585.1000 ;
      RECT 547.0500 582.1000 552.2000 585.1000 ;
      RECT 538.9000 582.1000 544.0500 585.1000 ;
      RECT 530.7500 582.1000 535.9000 585.1000 ;
      RECT 522.6000 582.1000 527.7500 585.1000 ;
      RECT 514.4500 582.1000 519.6000 585.1000 ;
      RECT 506.3000 582.1000 511.4500 585.1000 ;
      RECT 498.1500 582.1000 503.3000 585.1000 ;
      RECT 490.0000 582.1000 495.1500 585.1000 ;
      RECT 481.8500 582.1000 487.0000 585.1000 ;
      RECT 473.7000 582.1000 478.8500 585.1000 ;
      RECT 465.5500 582.1000 470.7000 585.1000 ;
      RECT 457.4000 582.1000 462.5500 585.1000 ;
      RECT 449.2500 582.1000 454.4000 585.1000 ;
      RECT 441.1000 582.1000 446.2500 585.1000 ;
      RECT 432.9500 582.1000 438.1000 585.1000 ;
      RECT 424.8000 582.1000 429.9500 585.1000 ;
      RECT 416.6500 582.1000 421.8000 585.1000 ;
      RECT 396.5000 582.1000 413.6500 585.1000 ;
      RECT 346.5000 582.1000 393.5000 585.1000 ;
      RECT 326.4650 582.1000 343.5000 585.1000 ;
      RECT 317.9500 582.1000 323.4650 585.1000 ;
      RECT 309.4350 582.1000 314.9500 585.1000 ;
      RECT 300.9200 582.1000 306.4350 585.1000 ;
      RECT 292.4050 582.1000 297.9200 585.1000 ;
      RECT 283.8900 582.1000 289.4050 585.1000 ;
      RECT 275.3750 582.1000 280.8900 585.1000 ;
      RECT 266.8600 582.1000 272.3750 585.1000 ;
      RECT 258.3450 582.1000 263.8600 585.1000 ;
      RECT 249.8300 582.1000 255.3450 585.1000 ;
      RECT 241.3150 582.1000 246.8300 585.1000 ;
      RECT 232.8000 582.1000 238.3150 585.1000 ;
      RECT 224.2850 582.1000 229.8000 585.1000 ;
      RECT 215.7700 582.1000 221.2850 585.1000 ;
      RECT 207.2550 582.1000 212.7700 585.1000 ;
      RECT 198.7400 582.1000 204.2550 585.1000 ;
      RECT 190.2250 582.1000 195.7400 585.1000 ;
      RECT 181.7100 582.1000 187.2250 585.1000 ;
      RECT 173.1950 582.1000 178.7100 585.1000 ;
      RECT 164.6800 582.1000 170.1950 585.1000 ;
      RECT 156.1650 582.1000 161.6800 585.1000 ;
      RECT 147.6500 582.1000 153.1650 585.1000 ;
      RECT 139.1350 582.1000 144.6500 585.1000 ;
      RECT 130.6200 582.1000 136.1350 585.1000 ;
      RECT 122.1050 582.1000 127.6200 585.1000 ;
      RECT 113.5900 582.1000 119.1050 585.1000 ;
      RECT 105.0750 582.1000 110.5900 585.1000 ;
      RECT 96.5600 582.1000 102.0750 585.1000 ;
      RECT 88.0450 582.1000 93.5600 585.1000 ;
      RECT 79.5300 582.1000 85.0450 585.1000 ;
      RECT 71.0150 582.1000 76.5300 585.1000 ;
      RECT 62.5000 582.1000 68.0150 585.1000 ;
      RECT 46.5000 582.1000 59.5000 585.1000 ;
      RECT 8.5000 582.1000 43.5000 585.1000 ;
      RECT 0.0000 582.1000 5.5000 585.1000 ;
      RECT 0.0000 580.7000 1120.0000 582.1000 ;
      RECT 1116.6000 580.1000 1120.0000 580.7000 ;
      RECT 0.0000 578.0050 1113.6000 580.7000 ;
      RECT 1118.5000 577.1000 1120.0000 580.1000 ;
      RECT 1114.5000 575.0050 1120.0000 577.1000 ;
      RECT 1076.5000 575.0050 1111.5000 578.0050 ;
      RECT 1060.5000 575.0050 1073.5000 578.0050 ;
      RECT 1052.3500 575.0050 1057.5000 578.0050 ;
      RECT 1044.2000 575.0050 1049.3500 578.0050 ;
      RECT 1036.0500 575.0050 1041.2000 578.0050 ;
      RECT 1027.9000 575.0050 1033.0500 578.0050 ;
      RECT 1019.7500 575.0050 1024.9000 578.0050 ;
      RECT 1011.6000 575.0050 1016.7500 578.0050 ;
      RECT 1003.4500 575.0050 1008.6000 578.0050 ;
      RECT 995.3000 575.0050 1000.4500 578.0050 ;
      RECT 987.1500 575.0050 992.3000 578.0050 ;
      RECT 979.0000 575.0050 984.1500 578.0050 ;
      RECT 970.8500 575.0050 976.0000 578.0050 ;
      RECT 962.7000 575.0050 967.8500 578.0050 ;
      RECT 954.5500 575.0050 959.7000 578.0050 ;
      RECT 946.4000 575.0050 951.5500 578.0050 ;
      RECT 938.2500 575.0050 943.4000 578.0050 ;
      RECT 930.1000 575.0050 935.2500 578.0050 ;
      RECT 921.9500 575.0050 927.1000 578.0050 ;
      RECT 913.8000 575.0050 918.9500 578.0050 ;
      RECT 905.6500 575.0050 910.8000 578.0050 ;
      RECT 897.5000 575.0050 902.6500 578.0050 ;
      RECT 889.3500 575.0050 894.5000 578.0050 ;
      RECT 881.2000 575.0050 886.3500 578.0050 ;
      RECT 873.0500 575.0050 878.2000 578.0050 ;
      RECT 864.9000 575.0050 870.0500 578.0050 ;
      RECT 856.7500 575.0050 861.9000 578.0050 ;
      RECT 848.6000 575.0050 853.7500 578.0050 ;
      RECT 840.4500 575.0050 845.6000 578.0050 ;
      RECT 832.3000 575.0050 837.4500 578.0050 ;
      RECT 824.1500 575.0050 829.3000 578.0050 ;
      RECT 816.0000 575.0050 821.1500 578.0050 ;
      RECT 807.8500 575.0050 813.0000 578.0050 ;
      RECT 799.7000 575.0050 804.8500 578.0050 ;
      RECT 791.5500 575.0050 796.7000 578.0050 ;
      RECT 783.4000 575.0050 788.5500 578.0050 ;
      RECT 775.2500 575.0050 780.4000 578.0050 ;
      RECT 767.1000 575.0050 772.2500 578.0050 ;
      RECT 758.9500 575.0050 764.1000 578.0050 ;
      RECT 750.8000 575.0050 755.9500 578.0050 ;
      RECT 742.6500 575.0050 747.8000 578.0050 ;
      RECT 734.5000 575.0050 739.6500 578.0050 ;
      RECT 726.3500 575.0050 731.5000 578.0050 ;
      RECT 718.2000 575.0050 723.3500 578.0050 ;
      RECT 710.0500 575.0050 715.2000 578.0050 ;
      RECT 701.9000 575.0050 707.0500 578.0050 ;
      RECT 693.7500 575.0050 698.9000 578.0050 ;
      RECT 685.6000 575.0050 690.7500 578.0050 ;
      RECT 677.4500 575.0050 682.6000 578.0050 ;
      RECT 669.3000 575.0050 674.4500 578.0050 ;
      RECT 661.1500 575.0050 666.3000 578.0050 ;
      RECT 653.0000 575.0050 658.1500 578.0050 ;
      RECT 644.8500 575.0050 650.0000 578.0050 ;
      RECT 636.7000 575.0050 641.8500 578.0050 ;
      RECT 628.5500 575.0050 633.7000 578.0050 ;
      RECT 620.4000 575.0050 625.5500 578.0050 ;
      RECT 612.2500 575.0050 617.4000 578.0050 ;
      RECT 604.1000 575.0050 609.2500 578.0050 ;
      RECT 595.9500 575.0050 601.1000 578.0050 ;
      RECT 587.8000 575.0050 592.9500 578.0050 ;
      RECT 579.6500 575.0050 584.8000 578.0050 ;
      RECT 571.5000 575.0050 576.6500 578.0050 ;
      RECT 563.3500 575.0050 568.5000 578.0050 ;
      RECT 555.2000 575.0050 560.3500 578.0050 ;
      RECT 547.0500 575.0050 552.2000 578.0050 ;
      RECT 538.9000 575.0050 544.0500 578.0050 ;
      RECT 530.7500 575.0050 535.9000 578.0050 ;
      RECT 522.6000 575.0050 527.7500 578.0050 ;
      RECT 514.4500 575.0050 519.6000 578.0050 ;
      RECT 506.3000 575.0050 511.4500 578.0050 ;
      RECT 498.1500 575.0050 503.3000 578.0050 ;
      RECT 490.0000 575.0050 495.1500 578.0050 ;
      RECT 481.8500 575.0050 487.0000 578.0050 ;
      RECT 473.7000 575.0050 478.8500 578.0050 ;
      RECT 465.5500 575.0050 470.7000 578.0050 ;
      RECT 457.4000 575.0050 462.5500 578.0050 ;
      RECT 449.2500 575.0050 454.4000 578.0050 ;
      RECT 441.1000 575.0050 446.2500 578.0050 ;
      RECT 432.9500 575.0050 438.1000 578.0050 ;
      RECT 424.8000 575.0050 429.9500 578.0050 ;
      RECT 416.6500 575.0050 421.8000 578.0050 ;
      RECT 396.5000 575.0050 413.6500 578.0050 ;
      RECT 346.5000 575.0050 393.5000 578.0050 ;
      RECT 326.4650 575.0050 343.5000 578.0050 ;
      RECT 317.9500 575.0050 323.4650 578.0050 ;
      RECT 309.4350 575.0050 314.9500 578.0050 ;
      RECT 300.9200 575.0050 306.4350 578.0050 ;
      RECT 292.4050 575.0050 297.9200 578.0050 ;
      RECT 283.8900 575.0050 289.4050 578.0050 ;
      RECT 275.3750 575.0050 280.8900 578.0050 ;
      RECT 266.8600 575.0050 272.3750 578.0050 ;
      RECT 258.3450 575.0050 263.8600 578.0050 ;
      RECT 249.8300 575.0050 255.3450 578.0050 ;
      RECT 241.3150 575.0050 246.8300 578.0050 ;
      RECT 232.8000 575.0050 238.3150 578.0050 ;
      RECT 224.2850 575.0050 229.8000 578.0050 ;
      RECT 215.7700 575.0050 221.2850 578.0050 ;
      RECT 207.2550 575.0050 212.7700 578.0050 ;
      RECT 198.7400 575.0050 204.2550 578.0050 ;
      RECT 190.2250 575.0050 195.7400 578.0050 ;
      RECT 181.7100 575.0050 187.2250 578.0050 ;
      RECT 173.1950 575.0050 178.7100 578.0050 ;
      RECT 164.6800 575.0050 170.1950 578.0050 ;
      RECT 156.1650 575.0050 161.6800 578.0050 ;
      RECT 147.6500 575.0050 153.1650 578.0050 ;
      RECT 139.1350 575.0050 144.6500 578.0050 ;
      RECT 130.6200 575.0050 136.1350 578.0050 ;
      RECT 122.1050 575.0050 127.6200 578.0050 ;
      RECT 113.5900 575.0050 119.1050 578.0050 ;
      RECT 105.0750 575.0050 110.5900 578.0050 ;
      RECT 96.5600 575.0050 102.0750 578.0050 ;
      RECT 88.0450 575.0050 93.5600 578.0050 ;
      RECT 79.5300 575.0050 85.0450 578.0050 ;
      RECT 71.0150 575.0050 76.5300 578.0050 ;
      RECT 62.5000 575.0050 68.0150 578.0050 ;
      RECT 46.5000 575.0050 59.5000 578.0050 ;
      RECT 8.5000 575.0050 43.5000 578.0050 ;
      RECT 0.0000 575.0050 5.5000 578.0050 ;
      RECT 0.0000 573.5000 1120.0000 575.0050 ;
      RECT 1116.6000 573.0050 1120.0000 573.5000 ;
      RECT 0.0000 570.9100 1113.6000 573.5000 ;
      RECT 1118.5000 570.0050 1120.0000 573.0050 ;
      RECT 1114.5000 567.9100 1120.0000 570.0050 ;
      RECT 1076.5000 567.9100 1111.5000 570.9100 ;
      RECT 1060.5000 567.9100 1073.5000 570.9100 ;
      RECT 1052.3500 567.9100 1057.5000 570.9100 ;
      RECT 1044.2000 567.9100 1049.3500 570.9100 ;
      RECT 1036.0500 567.9100 1041.2000 570.9100 ;
      RECT 1027.9000 567.9100 1033.0500 570.9100 ;
      RECT 1019.7500 567.9100 1024.9000 570.9100 ;
      RECT 1011.6000 567.9100 1016.7500 570.9100 ;
      RECT 1003.4500 567.9100 1008.6000 570.9100 ;
      RECT 995.3000 567.9100 1000.4500 570.9100 ;
      RECT 987.1500 567.9100 992.3000 570.9100 ;
      RECT 979.0000 567.9100 984.1500 570.9100 ;
      RECT 970.8500 567.9100 976.0000 570.9100 ;
      RECT 962.7000 567.9100 967.8500 570.9100 ;
      RECT 954.5500 567.9100 959.7000 570.9100 ;
      RECT 946.4000 567.9100 951.5500 570.9100 ;
      RECT 938.2500 567.9100 943.4000 570.9100 ;
      RECT 930.1000 567.9100 935.2500 570.9100 ;
      RECT 921.9500 567.9100 927.1000 570.9100 ;
      RECT 913.8000 567.9100 918.9500 570.9100 ;
      RECT 905.6500 567.9100 910.8000 570.9100 ;
      RECT 897.5000 567.9100 902.6500 570.9100 ;
      RECT 889.3500 567.9100 894.5000 570.9100 ;
      RECT 881.2000 567.9100 886.3500 570.9100 ;
      RECT 873.0500 567.9100 878.2000 570.9100 ;
      RECT 864.9000 567.9100 870.0500 570.9100 ;
      RECT 856.7500 567.9100 861.9000 570.9100 ;
      RECT 848.6000 567.9100 853.7500 570.9100 ;
      RECT 840.4500 567.9100 845.6000 570.9100 ;
      RECT 832.3000 567.9100 837.4500 570.9100 ;
      RECT 824.1500 567.9100 829.3000 570.9100 ;
      RECT 816.0000 567.9100 821.1500 570.9100 ;
      RECT 807.8500 567.9100 813.0000 570.9100 ;
      RECT 799.7000 567.9100 804.8500 570.9100 ;
      RECT 791.5500 567.9100 796.7000 570.9100 ;
      RECT 783.4000 567.9100 788.5500 570.9100 ;
      RECT 775.2500 567.9100 780.4000 570.9100 ;
      RECT 767.1000 567.9100 772.2500 570.9100 ;
      RECT 758.9500 567.9100 764.1000 570.9100 ;
      RECT 750.8000 567.9100 755.9500 570.9100 ;
      RECT 742.6500 567.9100 747.8000 570.9100 ;
      RECT 734.5000 567.9100 739.6500 570.9100 ;
      RECT 726.3500 567.9100 731.5000 570.9100 ;
      RECT 718.2000 567.9100 723.3500 570.9100 ;
      RECT 710.0500 567.9100 715.2000 570.9100 ;
      RECT 701.9000 567.9100 707.0500 570.9100 ;
      RECT 693.7500 567.9100 698.9000 570.9100 ;
      RECT 685.6000 567.9100 690.7500 570.9100 ;
      RECT 677.4500 567.9100 682.6000 570.9100 ;
      RECT 669.3000 567.9100 674.4500 570.9100 ;
      RECT 661.1500 567.9100 666.3000 570.9100 ;
      RECT 653.0000 567.9100 658.1500 570.9100 ;
      RECT 644.8500 567.9100 650.0000 570.9100 ;
      RECT 636.7000 567.9100 641.8500 570.9100 ;
      RECT 628.5500 567.9100 633.7000 570.9100 ;
      RECT 620.4000 567.9100 625.5500 570.9100 ;
      RECT 612.2500 567.9100 617.4000 570.9100 ;
      RECT 604.1000 567.9100 609.2500 570.9100 ;
      RECT 595.9500 567.9100 601.1000 570.9100 ;
      RECT 587.8000 567.9100 592.9500 570.9100 ;
      RECT 579.6500 567.9100 584.8000 570.9100 ;
      RECT 571.5000 567.9100 576.6500 570.9100 ;
      RECT 563.3500 567.9100 568.5000 570.9100 ;
      RECT 555.2000 567.9100 560.3500 570.9100 ;
      RECT 547.0500 567.9100 552.2000 570.9100 ;
      RECT 538.9000 567.9100 544.0500 570.9100 ;
      RECT 530.7500 567.9100 535.9000 570.9100 ;
      RECT 522.6000 567.9100 527.7500 570.9100 ;
      RECT 514.4500 567.9100 519.6000 570.9100 ;
      RECT 506.3000 567.9100 511.4500 570.9100 ;
      RECT 498.1500 567.9100 503.3000 570.9100 ;
      RECT 490.0000 567.9100 495.1500 570.9100 ;
      RECT 481.8500 567.9100 487.0000 570.9100 ;
      RECT 473.7000 567.9100 478.8500 570.9100 ;
      RECT 465.5500 567.9100 470.7000 570.9100 ;
      RECT 457.4000 567.9100 462.5500 570.9100 ;
      RECT 449.2500 567.9100 454.4000 570.9100 ;
      RECT 441.1000 567.9100 446.2500 570.9100 ;
      RECT 432.9500 567.9100 438.1000 570.9100 ;
      RECT 424.8000 567.9100 429.9500 570.9100 ;
      RECT 416.6500 567.9100 421.8000 570.9100 ;
      RECT 396.5000 567.9100 413.6500 570.9100 ;
      RECT 346.5000 567.9100 393.5000 570.9100 ;
      RECT 326.4650 567.9100 343.5000 570.9100 ;
      RECT 317.9500 567.9100 323.4650 570.9100 ;
      RECT 309.4350 567.9100 314.9500 570.9100 ;
      RECT 300.9200 567.9100 306.4350 570.9100 ;
      RECT 292.4050 567.9100 297.9200 570.9100 ;
      RECT 283.8900 567.9100 289.4050 570.9100 ;
      RECT 275.3750 567.9100 280.8900 570.9100 ;
      RECT 266.8600 567.9100 272.3750 570.9100 ;
      RECT 258.3450 567.9100 263.8600 570.9100 ;
      RECT 249.8300 567.9100 255.3450 570.9100 ;
      RECT 241.3150 567.9100 246.8300 570.9100 ;
      RECT 232.8000 567.9100 238.3150 570.9100 ;
      RECT 224.2850 567.9100 229.8000 570.9100 ;
      RECT 215.7700 567.9100 221.2850 570.9100 ;
      RECT 207.2550 567.9100 212.7700 570.9100 ;
      RECT 198.7400 567.9100 204.2550 570.9100 ;
      RECT 190.2250 567.9100 195.7400 570.9100 ;
      RECT 181.7100 567.9100 187.2250 570.9100 ;
      RECT 173.1950 567.9100 178.7100 570.9100 ;
      RECT 164.6800 567.9100 170.1950 570.9100 ;
      RECT 156.1650 567.9100 161.6800 570.9100 ;
      RECT 147.6500 567.9100 153.1650 570.9100 ;
      RECT 139.1350 567.9100 144.6500 570.9100 ;
      RECT 130.6200 567.9100 136.1350 570.9100 ;
      RECT 122.1050 567.9100 127.6200 570.9100 ;
      RECT 113.5900 567.9100 119.1050 570.9100 ;
      RECT 105.0750 567.9100 110.5900 570.9100 ;
      RECT 96.5600 567.9100 102.0750 570.9100 ;
      RECT 88.0450 567.9100 93.5600 570.9100 ;
      RECT 79.5300 567.9100 85.0450 570.9100 ;
      RECT 71.0150 567.9100 76.5300 570.9100 ;
      RECT 62.5000 567.9100 68.0150 570.9100 ;
      RECT 46.5000 567.9100 59.5000 570.9100 ;
      RECT 8.5000 567.9100 43.5000 570.9100 ;
      RECT 0.0000 567.9100 5.5000 570.9100 ;
      RECT 0.0000 566.5000 1120.0000 567.9100 ;
      RECT 1116.6000 565.9100 1120.0000 566.5000 ;
      RECT 0.0000 563.8150 1113.6000 566.5000 ;
      RECT 1118.5000 562.9100 1120.0000 565.9100 ;
      RECT 1114.5000 560.8150 1120.0000 562.9100 ;
      RECT 1076.5000 560.8150 1111.5000 563.8150 ;
      RECT 1060.5000 560.8150 1073.5000 563.8150 ;
      RECT 1052.3500 560.8150 1057.5000 563.8150 ;
      RECT 1044.2000 560.8150 1049.3500 563.8150 ;
      RECT 1036.0500 560.8150 1041.2000 563.8150 ;
      RECT 1027.9000 560.8150 1033.0500 563.8150 ;
      RECT 1019.7500 560.8150 1024.9000 563.8150 ;
      RECT 1011.6000 560.8150 1016.7500 563.8150 ;
      RECT 1003.4500 560.8150 1008.6000 563.8150 ;
      RECT 995.3000 560.8150 1000.4500 563.8150 ;
      RECT 987.1500 560.8150 992.3000 563.8150 ;
      RECT 979.0000 560.8150 984.1500 563.8150 ;
      RECT 970.8500 560.8150 976.0000 563.8150 ;
      RECT 962.7000 560.8150 967.8500 563.8150 ;
      RECT 954.5500 560.8150 959.7000 563.8150 ;
      RECT 946.4000 560.8150 951.5500 563.8150 ;
      RECT 938.2500 560.8150 943.4000 563.8150 ;
      RECT 930.1000 560.8150 935.2500 563.8150 ;
      RECT 921.9500 560.8150 927.1000 563.8150 ;
      RECT 913.8000 560.8150 918.9500 563.8150 ;
      RECT 905.6500 560.8150 910.8000 563.8150 ;
      RECT 897.5000 560.8150 902.6500 563.8150 ;
      RECT 889.3500 560.8150 894.5000 563.8150 ;
      RECT 881.2000 560.8150 886.3500 563.8150 ;
      RECT 873.0500 560.8150 878.2000 563.8150 ;
      RECT 864.9000 560.8150 870.0500 563.8150 ;
      RECT 856.7500 560.8150 861.9000 563.8150 ;
      RECT 848.6000 560.8150 853.7500 563.8150 ;
      RECT 840.4500 560.8150 845.6000 563.8150 ;
      RECT 832.3000 560.8150 837.4500 563.8150 ;
      RECT 824.1500 560.8150 829.3000 563.8150 ;
      RECT 816.0000 560.8150 821.1500 563.8150 ;
      RECT 807.8500 560.8150 813.0000 563.8150 ;
      RECT 799.7000 560.8150 804.8500 563.8150 ;
      RECT 791.5500 560.8150 796.7000 563.8150 ;
      RECT 783.4000 560.8150 788.5500 563.8150 ;
      RECT 775.2500 560.8150 780.4000 563.8150 ;
      RECT 767.1000 560.8150 772.2500 563.8150 ;
      RECT 758.9500 560.8150 764.1000 563.8150 ;
      RECT 750.8000 560.8150 755.9500 563.8150 ;
      RECT 742.6500 560.8150 747.8000 563.8150 ;
      RECT 734.5000 560.8150 739.6500 563.8150 ;
      RECT 726.3500 560.8150 731.5000 563.8150 ;
      RECT 718.2000 560.8150 723.3500 563.8150 ;
      RECT 710.0500 560.8150 715.2000 563.8150 ;
      RECT 701.9000 560.8150 707.0500 563.8150 ;
      RECT 693.7500 560.8150 698.9000 563.8150 ;
      RECT 685.6000 560.8150 690.7500 563.8150 ;
      RECT 677.4500 560.8150 682.6000 563.8150 ;
      RECT 669.3000 560.8150 674.4500 563.8150 ;
      RECT 661.1500 560.8150 666.3000 563.8150 ;
      RECT 653.0000 560.8150 658.1500 563.8150 ;
      RECT 644.8500 560.8150 650.0000 563.8150 ;
      RECT 636.7000 560.8150 641.8500 563.8150 ;
      RECT 628.5500 560.8150 633.7000 563.8150 ;
      RECT 620.4000 560.8150 625.5500 563.8150 ;
      RECT 612.2500 560.8150 617.4000 563.8150 ;
      RECT 604.1000 560.8150 609.2500 563.8150 ;
      RECT 595.9500 560.8150 601.1000 563.8150 ;
      RECT 587.8000 560.8150 592.9500 563.8150 ;
      RECT 579.6500 560.8150 584.8000 563.8150 ;
      RECT 571.5000 560.8150 576.6500 563.8150 ;
      RECT 563.3500 560.8150 568.5000 563.8150 ;
      RECT 555.2000 560.8150 560.3500 563.8150 ;
      RECT 547.0500 560.8150 552.2000 563.8150 ;
      RECT 538.9000 560.8150 544.0500 563.8150 ;
      RECT 530.7500 560.8150 535.9000 563.8150 ;
      RECT 522.6000 560.8150 527.7500 563.8150 ;
      RECT 514.4500 560.8150 519.6000 563.8150 ;
      RECT 506.3000 560.8150 511.4500 563.8150 ;
      RECT 498.1500 560.8150 503.3000 563.8150 ;
      RECT 490.0000 560.8150 495.1500 563.8150 ;
      RECT 481.8500 560.8150 487.0000 563.8150 ;
      RECT 473.7000 560.8150 478.8500 563.8150 ;
      RECT 465.5500 560.8150 470.7000 563.8150 ;
      RECT 457.4000 560.8150 462.5500 563.8150 ;
      RECT 449.2500 560.8150 454.4000 563.8150 ;
      RECT 441.1000 560.8150 446.2500 563.8150 ;
      RECT 432.9500 560.8150 438.1000 563.8150 ;
      RECT 424.8000 560.8150 429.9500 563.8150 ;
      RECT 416.6500 560.8150 421.8000 563.8150 ;
      RECT 396.5000 560.8150 413.6500 563.8150 ;
      RECT 346.5000 560.8150 393.5000 563.8150 ;
      RECT 326.4650 560.8150 343.5000 563.8150 ;
      RECT 317.9500 560.8150 323.4650 563.8150 ;
      RECT 309.4350 560.8150 314.9500 563.8150 ;
      RECT 300.9200 560.8150 306.4350 563.8150 ;
      RECT 292.4050 560.8150 297.9200 563.8150 ;
      RECT 283.8900 560.8150 289.4050 563.8150 ;
      RECT 275.3750 560.8150 280.8900 563.8150 ;
      RECT 266.8600 560.8150 272.3750 563.8150 ;
      RECT 258.3450 560.8150 263.8600 563.8150 ;
      RECT 249.8300 560.8150 255.3450 563.8150 ;
      RECT 241.3150 560.8150 246.8300 563.8150 ;
      RECT 232.8000 560.8150 238.3150 563.8150 ;
      RECT 224.2850 560.8150 229.8000 563.8150 ;
      RECT 215.7700 560.8150 221.2850 563.8150 ;
      RECT 207.2550 560.8150 212.7700 563.8150 ;
      RECT 198.7400 560.8150 204.2550 563.8150 ;
      RECT 190.2250 560.8150 195.7400 563.8150 ;
      RECT 181.7100 560.8150 187.2250 563.8150 ;
      RECT 173.1950 560.8150 178.7100 563.8150 ;
      RECT 164.6800 560.8150 170.1950 563.8150 ;
      RECT 156.1650 560.8150 161.6800 563.8150 ;
      RECT 147.6500 560.8150 153.1650 563.8150 ;
      RECT 139.1350 560.8150 144.6500 563.8150 ;
      RECT 130.6200 560.8150 136.1350 563.8150 ;
      RECT 122.1050 560.8150 127.6200 563.8150 ;
      RECT 113.5900 560.8150 119.1050 563.8150 ;
      RECT 105.0750 560.8150 110.5900 563.8150 ;
      RECT 96.5600 560.8150 102.0750 563.8150 ;
      RECT 88.0450 560.8150 93.5600 563.8150 ;
      RECT 79.5300 560.8150 85.0450 563.8150 ;
      RECT 71.0150 560.8150 76.5300 563.8150 ;
      RECT 62.5000 560.8150 68.0150 563.8150 ;
      RECT 46.5000 560.8150 59.5000 563.8150 ;
      RECT 8.5000 560.8150 43.5000 563.8150 ;
      RECT 0.0000 560.8150 5.5000 563.8150 ;
      RECT 0.0000 559.3000 1120.0000 560.8150 ;
      RECT 1116.6000 558.8150 1120.0000 559.3000 ;
      RECT 0.0000 556.7200 1113.6000 559.3000 ;
      RECT 1118.5000 555.8150 1120.0000 558.8150 ;
      RECT 1114.5000 553.7200 1120.0000 555.8150 ;
      RECT 1076.5000 553.7200 1111.5000 556.7200 ;
      RECT 1060.5000 553.7200 1073.5000 556.7200 ;
      RECT 1052.3500 553.7200 1057.5000 556.7200 ;
      RECT 1044.2000 553.7200 1049.3500 556.7200 ;
      RECT 1036.0500 553.7200 1041.2000 556.7200 ;
      RECT 1027.9000 553.7200 1033.0500 556.7200 ;
      RECT 1019.7500 553.7200 1024.9000 556.7200 ;
      RECT 1011.6000 553.7200 1016.7500 556.7200 ;
      RECT 1003.4500 553.7200 1008.6000 556.7200 ;
      RECT 995.3000 553.7200 1000.4500 556.7200 ;
      RECT 987.1500 553.7200 992.3000 556.7200 ;
      RECT 979.0000 553.7200 984.1500 556.7200 ;
      RECT 970.8500 553.7200 976.0000 556.7200 ;
      RECT 962.7000 553.7200 967.8500 556.7200 ;
      RECT 954.5500 553.7200 959.7000 556.7200 ;
      RECT 946.4000 553.7200 951.5500 556.7200 ;
      RECT 938.2500 553.7200 943.4000 556.7200 ;
      RECT 930.1000 553.7200 935.2500 556.7200 ;
      RECT 921.9500 553.7200 927.1000 556.7200 ;
      RECT 913.8000 553.7200 918.9500 556.7200 ;
      RECT 905.6500 553.7200 910.8000 556.7200 ;
      RECT 897.5000 553.7200 902.6500 556.7200 ;
      RECT 889.3500 553.7200 894.5000 556.7200 ;
      RECT 881.2000 553.7200 886.3500 556.7200 ;
      RECT 873.0500 553.7200 878.2000 556.7200 ;
      RECT 864.9000 553.7200 870.0500 556.7200 ;
      RECT 856.7500 553.7200 861.9000 556.7200 ;
      RECT 848.6000 553.7200 853.7500 556.7200 ;
      RECT 840.4500 553.7200 845.6000 556.7200 ;
      RECT 832.3000 553.7200 837.4500 556.7200 ;
      RECT 824.1500 553.7200 829.3000 556.7200 ;
      RECT 816.0000 553.7200 821.1500 556.7200 ;
      RECT 807.8500 553.7200 813.0000 556.7200 ;
      RECT 799.7000 553.7200 804.8500 556.7200 ;
      RECT 791.5500 553.7200 796.7000 556.7200 ;
      RECT 783.4000 553.7200 788.5500 556.7200 ;
      RECT 775.2500 553.7200 780.4000 556.7200 ;
      RECT 767.1000 553.7200 772.2500 556.7200 ;
      RECT 758.9500 553.7200 764.1000 556.7200 ;
      RECT 750.8000 553.7200 755.9500 556.7200 ;
      RECT 742.6500 553.7200 747.8000 556.7200 ;
      RECT 734.5000 553.7200 739.6500 556.7200 ;
      RECT 726.3500 553.7200 731.5000 556.7200 ;
      RECT 718.2000 553.7200 723.3500 556.7200 ;
      RECT 710.0500 553.7200 715.2000 556.7200 ;
      RECT 701.9000 553.7200 707.0500 556.7200 ;
      RECT 693.7500 553.7200 698.9000 556.7200 ;
      RECT 685.6000 553.7200 690.7500 556.7200 ;
      RECT 677.4500 553.7200 682.6000 556.7200 ;
      RECT 669.3000 553.7200 674.4500 556.7200 ;
      RECT 661.1500 553.7200 666.3000 556.7200 ;
      RECT 653.0000 553.7200 658.1500 556.7200 ;
      RECT 644.8500 553.7200 650.0000 556.7200 ;
      RECT 636.7000 553.7200 641.8500 556.7200 ;
      RECT 628.5500 553.7200 633.7000 556.7200 ;
      RECT 620.4000 553.7200 625.5500 556.7200 ;
      RECT 612.2500 553.7200 617.4000 556.7200 ;
      RECT 604.1000 553.7200 609.2500 556.7200 ;
      RECT 595.9500 553.7200 601.1000 556.7200 ;
      RECT 587.8000 553.7200 592.9500 556.7200 ;
      RECT 579.6500 553.7200 584.8000 556.7200 ;
      RECT 571.5000 553.7200 576.6500 556.7200 ;
      RECT 563.3500 553.7200 568.5000 556.7200 ;
      RECT 555.2000 553.7200 560.3500 556.7200 ;
      RECT 547.0500 553.7200 552.2000 556.7200 ;
      RECT 538.9000 553.7200 544.0500 556.7200 ;
      RECT 530.7500 553.7200 535.9000 556.7200 ;
      RECT 522.6000 553.7200 527.7500 556.7200 ;
      RECT 514.4500 553.7200 519.6000 556.7200 ;
      RECT 506.3000 553.7200 511.4500 556.7200 ;
      RECT 498.1500 553.7200 503.3000 556.7200 ;
      RECT 490.0000 553.7200 495.1500 556.7200 ;
      RECT 481.8500 553.7200 487.0000 556.7200 ;
      RECT 473.7000 553.7200 478.8500 556.7200 ;
      RECT 465.5500 553.7200 470.7000 556.7200 ;
      RECT 457.4000 553.7200 462.5500 556.7200 ;
      RECT 449.2500 553.7200 454.4000 556.7200 ;
      RECT 441.1000 553.7200 446.2500 556.7200 ;
      RECT 432.9500 553.7200 438.1000 556.7200 ;
      RECT 424.8000 553.7200 429.9500 556.7200 ;
      RECT 416.6500 553.7200 421.8000 556.7200 ;
      RECT 396.5000 553.7200 413.6500 556.7200 ;
      RECT 346.5000 553.7200 393.5000 556.7200 ;
      RECT 326.4650 553.7200 343.5000 556.7200 ;
      RECT 317.9500 553.7200 323.4650 556.7200 ;
      RECT 309.4350 553.7200 314.9500 556.7200 ;
      RECT 300.9200 553.7200 306.4350 556.7200 ;
      RECT 292.4050 553.7200 297.9200 556.7200 ;
      RECT 283.8900 553.7200 289.4050 556.7200 ;
      RECT 275.3750 553.7200 280.8900 556.7200 ;
      RECT 266.8600 553.7200 272.3750 556.7200 ;
      RECT 258.3450 553.7200 263.8600 556.7200 ;
      RECT 249.8300 553.7200 255.3450 556.7200 ;
      RECT 241.3150 553.7200 246.8300 556.7200 ;
      RECT 232.8000 553.7200 238.3150 556.7200 ;
      RECT 224.2850 553.7200 229.8000 556.7200 ;
      RECT 215.7700 553.7200 221.2850 556.7200 ;
      RECT 207.2550 553.7200 212.7700 556.7200 ;
      RECT 198.7400 553.7200 204.2550 556.7200 ;
      RECT 190.2250 553.7200 195.7400 556.7200 ;
      RECT 181.7100 553.7200 187.2250 556.7200 ;
      RECT 173.1950 553.7200 178.7100 556.7200 ;
      RECT 164.6800 553.7200 170.1950 556.7200 ;
      RECT 156.1650 553.7200 161.6800 556.7200 ;
      RECT 147.6500 553.7200 153.1650 556.7200 ;
      RECT 139.1350 553.7200 144.6500 556.7200 ;
      RECT 130.6200 553.7200 136.1350 556.7200 ;
      RECT 122.1050 553.7200 127.6200 556.7200 ;
      RECT 113.5900 553.7200 119.1050 556.7200 ;
      RECT 105.0750 553.7200 110.5900 556.7200 ;
      RECT 96.5600 553.7200 102.0750 556.7200 ;
      RECT 88.0450 553.7200 93.5600 556.7200 ;
      RECT 79.5300 553.7200 85.0450 556.7200 ;
      RECT 71.0150 553.7200 76.5300 556.7200 ;
      RECT 62.5000 553.7200 68.0150 556.7200 ;
      RECT 46.5000 553.7200 59.5000 556.7200 ;
      RECT 8.5000 553.7200 43.5000 556.7200 ;
      RECT 0.0000 553.7200 5.5000 556.7200 ;
      RECT 0.0000 552.3000 1120.0000 553.7200 ;
      RECT 1116.6000 551.7200 1120.0000 552.3000 ;
      RECT 0.0000 549.6250 1113.6000 552.3000 ;
      RECT 1118.5000 548.7200 1120.0000 551.7200 ;
      RECT 1114.5000 546.6250 1120.0000 548.7200 ;
      RECT 1076.5000 546.6250 1111.5000 549.6250 ;
      RECT 1060.5000 546.6250 1073.5000 549.6250 ;
      RECT 1052.3500 546.6250 1057.5000 549.6250 ;
      RECT 1044.2000 546.6250 1049.3500 549.6250 ;
      RECT 1036.0500 546.6250 1041.2000 549.6250 ;
      RECT 1027.9000 546.6250 1033.0500 549.6250 ;
      RECT 1019.7500 546.6250 1024.9000 549.6250 ;
      RECT 1011.6000 546.6250 1016.7500 549.6250 ;
      RECT 1003.4500 546.6250 1008.6000 549.6250 ;
      RECT 995.3000 546.6250 1000.4500 549.6250 ;
      RECT 987.1500 546.6250 992.3000 549.6250 ;
      RECT 979.0000 546.6250 984.1500 549.6250 ;
      RECT 970.8500 546.6250 976.0000 549.6250 ;
      RECT 962.7000 546.6250 967.8500 549.6250 ;
      RECT 954.5500 546.6250 959.7000 549.6250 ;
      RECT 946.4000 546.6250 951.5500 549.6250 ;
      RECT 938.2500 546.6250 943.4000 549.6250 ;
      RECT 930.1000 546.6250 935.2500 549.6250 ;
      RECT 921.9500 546.6250 927.1000 549.6250 ;
      RECT 913.8000 546.6250 918.9500 549.6250 ;
      RECT 905.6500 546.6250 910.8000 549.6250 ;
      RECT 897.5000 546.6250 902.6500 549.6250 ;
      RECT 889.3500 546.6250 894.5000 549.6250 ;
      RECT 881.2000 546.6250 886.3500 549.6250 ;
      RECT 873.0500 546.6250 878.2000 549.6250 ;
      RECT 864.9000 546.6250 870.0500 549.6250 ;
      RECT 856.7500 546.6250 861.9000 549.6250 ;
      RECT 848.6000 546.6250 853.7500 549.6250 ;
      RECT 840.4500 546.6250 845.6000 549.6250 ;
      RECT 832.3000 546.6250 837.4500 549.6250 ;
      RECT 824.1500 546.6250 829.3000 549.6250 ;
      RECT 816.0000 546.6250 821.1500 549.6250 ;
      RECT 807.8500 546.6250 813.0000 549.6250 ;
      RECT 799.7000 546.6250 804.8500 549.6250 ;
      RECT 791.5500 546.6250 796.7000 549.6250 ;
      RECT 783.4000 546.6250 788.5500 549.6250 ;
      RECT 775.2500 546.6250 780.4000 549.6250 ;
      RECT 767.1000 546.6250 772.2500 549.6250 ;
      RECT 758.9500 546.6250 764.1000 549.6250 ;
      RECT 750.8000 546.6250 755.9500 549.6250 ;
      RECT 742.6500 546.6250 747.8000 549.6250 ;
      RECT 734.5000 546.6250 739.6500 549.6250 ;
      RECT 726.3500 546.6250 731.5000 549.6250 ;
      RECT 718.2000 546.6250 723.3500 549.6250 ;
      RECT 710.0500 546.6250 715.2000 549.6250 ;
      RECT 701.9000 546.6250 707.0500 549.6250 ;
      RECT 693.7500 546.6250 698.9000 549.6250 ;
      RECT 685.6000 546.6250 690.7500 549.6250 ;
      RECT 677.4500 546.6250 682.6000 549.6250 ;
      RECT 669.3000 546.6250 674.4500 549.6250 ;
      RECT 661.1500 546.6250 666.3000 549.6250 ;
      RECT 653.0000 546.6250 658.1500 549.6250 ;
      RECT 644.8500 546.6250 650.0000 549.6250 ;
      RECT 636.7000 546.6250 641.8500 549.6250 ;
      RECT 628.5500 546.6250 633.7000 549.6250 ;
      RECT 620.4000 546.6250 625.5500 549.6250 ;
      RECT 612.2500 546.6250 617.4000 549.6250 ;
      RECT 604.1000 546.6250 609.2500 549.6250 ;
      RECT 595.9500 546.6250 601.1000 549.6250 ;
      RECT 587.8000 546.6250 592.9500 549.6250 ;
      RECT 579.6500 546.6250 584.8000 549.6250 ;
      RECT 571.5000 546.6250 576.6500 549.6250 ;
      RECT 563.3500 546.6250 568.5000 549.6250 ;
      RECT 555.2000 546.6250 560.3500 549.6250 ;
      RECT 547.0500 546.6250 552.2000 549.6250 ;
      RECT 538.9000 546.6250 544.0500 549.6250 ;
      RECT 530.7500 546.6250 535.9000 549.6250 ;
      RECT 522.6000 546.6250 527.7500 549.6250 ;
      RECT 514.4500 546.6250 519.6000 549.6250 ;
      RECT 506.3000 546.6250 511.4500 549.6250 ;
      RECT 498.1500 546.6250 503.3000 549.6250 ;
      RECT 490.0000 546.6250 495.1500 549.6250 ;
      RECT 481.8500 546.6250 487.0000 549.6250 ;
      RECT 473.7000 546.6250 478.8500 549.6250 ;
      RECT 465.5500 546.6250 470.7000 549.6250 ;
      RECT 457.4000 546.6250 462.5500 549.6250 ;
      RECT 449.2500 546.6250 454.4000 549.6250 ;
      RECT 441.1000 546.6250 446.2500 549.6250 ;
      RECT 432.9500 546.6250 438.1000 549.6250 ;
      RECT 424.8000 546.6250 429.9500 549.6250 ;
      RECT 416.6500 546.6250 421.8000 549.6250 ;
      RECT 396.5000 546.6250 413.6500 549.6250 ;
      RECT 346.5000 546.6250 393.5000 549.6250 ;
      RECT 326.4650 546.6250 343.5000 549.6250 ;
      RECT 317.9500 546.6250 323.4650 549.6250 ;
      RECT 309.4350 546.6250 314.9500 549.6250 ;
      RECT 300.9200 546.6250 306.4350 549.6250 ;
      RECT 292.4050 546.6250 297.9200 549.6250 ;
      RECT 283.8900 546.6250 289.4050 549.6250 ;
      RECT 275.3750 546.6250 280.8900 549.6250 ;
      RECT 266.8600 546.6250 272.3750 549.6250 ;
      RECT 258.3450 546.6250 263.8600 549.6250 ;
      RECT 249.8300 546.6250 255.3450 549.6250 ;
      RECT 241.3150 546.6250 246.8300 549.6250 ;
      RECT 232.8000 546.6250 238.3150 549.6250 ;
      RECT 224.2850 546.6250 229.8000 549.6250 ;
      RECT 215.7700 546.6250 221.2850 549.6250 ;
      RECT 207.2550 546.6250 212.7700 549.6250 ;
      RECT 198.7400 546.6250 204.2550 549.6250 ;
      RECT 190.2250 546.6250 195.7400 549.6250 ;
      RECT 181.7100 546.6250 187.2250 549.6250 ;
      RECT 173.1950 546.6250 178.7100 549.6250 ;
      RECT 164.6800 546.6250 170.1950 549.6250 ;
      RECT 156.1650 546.6250 161.6800 549.6250 ;
      RECT 147.6500 546.6250 153.1650 549.6250 ;
      RECT 139.1350 546.6250 144.6500 549.6250 ;
      RECT 130.6200 546.6250 136.1350 549.6250 ;
      RECT 122.1050 546.6250 127.6200 549.6250 ;
      RECT 113.5900 546.6250 119.1050 549.6250 ;
      RECT 105.0750 546.6250 110.5900 549.6250 ;
      RECT 96.5600 546.6250 102.0750 549.6250 ;
      RECT 88.0450 546.6250 93.5600 549.6250 ;
      RECT 79.5300 546.6250 85.0450 549.6250 ;
      RECT 71.0150 546.6250 76.5300 549.6250 ;
      RECT 62.5000 546.6250 68.0150 549.6250 ;
      RECT 46.5000 546.6250 59.5000 549.6250 ;
      RECT 8.5000 546.6250 43.5000 549.6250 ;
      RECT 0.0000 546.6250 5.5000 549.6250 ;
      RECT 0.0000 545.1000 1120.0000 546.6250 ;
      RECT 1116.6000 544.6250 1120.0000 545.1000 ;
      RECT 0.0000 542.5300 1113.6000 545.1000 ;
      RECT 1118.5000 541.6250 1120.0000 544.6250 ;
      RECT 1114.5000 539.5300 1120.0000 541.6250 ;
      RECT 1076.5000 539.5300 1111.5000 542.5300 ;
      RECT 1060.5000 539.5300 1073.5000 542.5300 ;
      RECT 1052.3500 539.5300 1057.5000 542.5300 ;
      RECT 1044.2000 539.5300 1049.3500 542.5300 ;
      RECT 1036.0500 539.5300 1041.2000 542.5300 ;
      RECT 1027.9000 539.5300 1033.0500 542.5300 ;
      RECT 1019.7500 539.5300 1024.9000 542.5300 ;
      RECT 1011.6000 539.5300 1016.7500 542.5300 ;
      RECT 1003.4500 539.5300 1008.6000 542.5300 ;
      RECT 995.3000 539.5300 1000.4500 542.5300 ;
      RECT 987.1500 539.5300 992.3000 542.5300 ;
      RECT 979.0000 539.5300 984.1500 542.5300 ;
      RECT 970.8500 539.5300 976.0000 542.5300 ;
      RECT 962.7000 539.5300 967.8500 542.5300 ;
      RECT 954.5500 539.5300 959.7000 542.5300 ;
      RECT 946.4000 539.5300 951.5500 542.5300 ;
      RECT 938.2500 539.5300 943.4000 542.5300 ;
      RECT 930.1000 539.5300 935.2500 542.5300 ;
      RECT 921.9500 539.5300 927.1000 542.5300 ;
      RECT 913.8000 539.5300 918.9500 542.5300 ;
      RECT 905.6500 539.5300 910.8000 542.5300 ;
      RECT 897.5000 539.5300 902.6500 542.5300 ;
      RECT 889.3500 539.5300 894.5000 542.5300 ;
      RECT 881.2000 539.5300 886.3500 542.5300 ;
      RECT 873.0500 539.5300 878.2000 542.5300 ;
      RECT 864.9000 539.5300 870.0500 542.5300 ;
      RECT 856.7500 539.5300 861.9000 542.5300 ;
      RECT 848.6000 539.5300 853.7500 542.5300 ;
      RECT 840.4500 539.5300 845.6000 542.5300 ;
      RECT 832.3000 539.5300 837.4500 542.5300 ;
      RECT 824.1500 539.5300 829.3000 542.5300 ;
      RECT 816.0000 539.5300 821.1500 542.5300 ;
      RECT 807.8500 539.5300 813.0000 542.5300 ;
      RECT 799.7000 539.5300 804.8500 542.5300 ;
      RECT 791.5500 539.5300 796.7000 542.5300 ;
      RECT 783.4000 539.5300 788.5500 542.5300 ;
      RECT 775.2500 539.5300 780.4000 542.5300 ;
      RECT 767.1000 539.5300 772.2500 542.5300 ;
      RECT 758.9500 539.5300 764.1000 542.5300 ;
      RECT 750.8000 539.5300 755.9500 542.5300 ;
      RECT 742.6500 539.5300 747.8000 542.5300 ;
      RECT 734.5000 539.5300 739.6500 542.5300 ;
      RECT 726.3500 539.5300 731.5000 542.5300 ;
      RECT 718.2000 539.5300 723.3500 542.5300 ;
      RECT 710.0500 539.5300 715.2000 542.5300 ;
      RECT 701.9000 539.5300 707.0500 542.5300 ;
      RECT 693.7500 539.5300 698.9000 542.5300 ;
      RECT 685.6000 539.5300 690.7500 542.5300 ;
      RECT 677.4500 539.5300 682.6000 542.5300 ;
      RECT 669.3000 539.5300 674.4500 542.5300 ;
      RECT 661.1500 539.5300 666.3000 542.5300 ;
      RECT 653.0000 539.5300 658.1500 542.5300 ;
      RECT 644.8500 539.5300 650.0000 542.5300 ;
      RECT 636.7000 539.5300 641.8500 542.5300 ;
      RECT 628.5500 539.5300 633.7000 542.5300 ;
      RECT 620.4000 539.5300 625.5500 542.5300 ;
      RECT 612.2500 539.5300 617.4000 542.5300 ;
      RECT 604.1000 539.5300 609.2500 542.5300 ;
      RECT 595.9500 539.5300 601.1000 542.5300 ;
      RECT 587.8000 539.5300 592.9500 542.5300 ;
      RECT 579.6500 539.5300 584.8000 542.5300 ;
      RECT 571.5000 539.5300 576.6500 542.5300 ;
      RECT 563.3500 539.5300 568.5000 542.5300 ;
      RECT 555.2000 539.5300 560.3500 542.5300 ;
      RECT 547.0500 539.5300 552.2000 542.5300 ;
      RECT 538.9000 539.5300 544.0500 542.5300 ;
      RECT 530.7500 539.5300 535.9000 542.5300 ;
      RECT 522.6000 539.5300 527.7500 542.5300 ;
      RECT 514.4500 539.5300 519.6000 542.5300 ;
      RECT 506.3000 539.5300 511.4500 542.5300 ;
      RECT 498.1500 539.5300 503.3000 542.5300 ;
      RECT 490.0000 539.5300 495.1500 542.5300 ;
      RECT 481.8500 539.5300 487.0000 542.5300 ;
      RECT 473.7000 539.5300 478.8500 542.5300 ;
      RECT 465.5500 539.5300 470.7000 542.5300 ;
      RECT 457.4000 539.5300 462.5500 542.5300 ;
      RECT 449.2500 539.5300 454.4000 542.5300 ;
      RECT 441.1000 539.5300 446.2500 542.5300 ;
      RECT 432.9500 539.5300 438.1000 542.5300 ;
      RECT 424.8000 539.5300 429.9500 542.5300 ;
      RECT 416.6500 539.5300 421.8000 542.5300 ;
      RECT 396.5000 539.5300 413.6500 542.5300 ;
      RECT 346.5000 539.5300 393.5000 542.5300 ;
      RECT 326.4650 539.5300 343.5000 542.5300 ;
      RECT 317.9500 539.5300 323.4650 542.5300 ;
      RECT 309.4350 539.5300 314.9500 542.5300 ;
      RECT 300.9200 539.5300 306.4350 542.5300 ;
      RECT 292.4050 539.5300 297.9200 542.5300 ;
      RECT 283.8900 539.5300 289.4050 542.5300 ;
      RECT 275.3750 539.5300 280.8900 542.5300 ;
      RECT 266.8600 539.5300 272.3750 542.5300 ;
      RECT 258.3450 539.5300 263.8600 542.5300 ;
      RECT 249.8300 539.5300 255.3450 542.5300 ;
      RECT 241.3150 539.5300 246.8300 542.5300 ;
      RECT 232.8000 539.5300 238.3150 542.5300 ;
      RECT 224.2850 539.5300 229.8000 542.5300 ;
      RECT 215.7700 539.5300 221.2850 542.5300 ;
      RECT 207.2550 539.5300 212.7700 542.5300 ;
      RECT 198.7400 539.5300 204.2550 542.5300 ;
      RECT 190.2250 539.5300 195.7400 542.5300 ;
      RECT 181.7100 539.5300 187.2250 542.5300 ;
      RECT 173.1950 539.5300 178.7100 542.5300 ;
      RECT 164.6800 539.5300 170.1950 542.5300 ;
      RECT 156.1650 539.5300 161.6800 542.5300 ;
      RECT 147.6500 539.5300 153.1650 542.5300 ;
      RECT 139.1350 539.5300 144.6500 542.5300 ;
      RECT 130.6200 539.5300 136.1350 542.5300 ;
      RECT 122.1050 539.5300 127.6200 542.5300 ;
      RECT 113.5900 539.5300 119.1050 542.5300 ;
      RECT 105.0750 539.5300 110.5900 542.5300 ;
      RECT 96.5600 539.5300 102.0750 542.5300 ;
      RECT 88.0450 539.5300 93.5600 542.5300 ;
      RECT 79.5300 539.5300 85.0450 542.5300 ;
      RECT 71.0150 539.5300 76.5300 542.5300 ;
      RECT 62.5000 539.5300 68.0150 542.5300 ;
      RECT 46.5000 539.5300 59.5000 542.5300 ;
      RECT 8.5000 539.5300 43.5000 542.5300 ;
      RECT 0.0000 539.5300 5.5000 542.5300 ;
      RECT 0.0000 538.1000 1120.0000 539.5300 ;
      RECT 1116.6000 537.5300 1120.0000 538.1000 ;
      RECT 0.0000 535.4350 1113.6000 538.1000 ;
      RECT 1118.5000 534.5300 1120.0000 537.5300 ;
      RECT 1114.5000 532.4350 1120.0000 534.5300 ;
      RECT 1076.5000 532.4350 1111.5000 535.4350 ;
      RECT 1060.5000 532.4350 1073.5000 535.4350 ;
      RECT 1052.3500 532.4350 1057.5000 535.4350 ;
      RECT 1044.2000 532.4350 1049.3500 535.4350 ;
      RECT 1036.0500 532.4350 1041.2000 535.4350 ;
      RECT 1027.9000 532.4350 1033.0500 535.4350 ;
      RECT 1019.7500 532.4350 1024.9000 535.4350 ;
      RECT 1011.6000 532.4350 1016.7500 535.4350 ;
      RECT 1003.4500 532.4350 1008.6000 535.4350 ;
      RECT 995.3000 532.4350 1000.4500 535.4350 ;
      RECT 987.1500 532.4350 992.3000 535.4350 ;
      RECT 979.0000 532.4350 984.1500 535.4350 ;
      RECT 970.8500 532.4350 976.0000 535.4350 ;
      RECT 962.7000 532.4350 967.8500 535.4350 ;
      RECT 954.5500 532.4350 959.7000 535.4350 ;
      RECT 946.4000 532.4350 951.5500 535.4350 ;
      RECT 938.2500 532.4350 943.4000 535.4350 ;
      RECT 930.1000 532.4350 935.2500 535.4350 ;
      RECT 921.9500 532.4350 927.1000 535.4350 ;
      RECT 913.8000 532.4350 918.9500 535.4350 ;
      RECT 905.6500 532.4350 910.8000 535.4350 ;
      RECT 897.5000 532.4350 902.6500 535.4350 ;
      RECT 889.3500 532.4350 894.5000 535.4350 ;
      RECT 881.2000 532.4350 886.3500 535.4350 ;
      RECT 873.0500 532.4350 878.2000 535.4350 ;
      RECT 864.9000 532.4350 870.0500 535.4350 ;
      RECT 856.7500 532.4350 861.9000 535.4350 ;
      RECT 848.6000 532.4350 853.7500 535.4350 ;
      RECT 840.4500 532.4350 845.6000 535.4350 ;
      RECT 832.3000 532.4350 837.4500 535.4350 ;
      RECT 824.1500 532.4350 829.3000 535.4350 ;
      RECT 816.0000 532.4350 821.1500 535.4350 ;
      RECT 807.8500 532.4350 813.0000 535.4350 ;
      RECT 799.7000 532.4350 804.8500 535.4350 ;
      RECT 791.5500 532.4350 796.7000 535.4350 ;
      RECT 783.4000 532.4350 788.5500 535.4350 ;
      RECT 775.2500 532.4350 780.4000 535.4350 ;
      RECT 767.1000 532.4350 772.2500 535.4350 ;
      RECT 758.9500 532.4350 764.1000 535.4350 ;
      RECT 750.8000 532.4350 755.9500 535.4350 ;
      RECT 742.6500 532.4350 747.8000 535.4350 ;
      RECT 734.5000 532.4350 739.6500 535.4350 ;
      RECT 726.3500 532.4350 731.5000 535.4350 ;
      RECT 718.2000 532.4350 723.3500 535.4350 ;
      RECT 710.0500 532.4350 715.2000 535.4350 ;
      RECT 701.9000 532.4350 707.0500 535.4350 ;
      RECT 693.7500 532.4350 698.9000 535.4350 ;
      RECT 685.6000 532.4350 690.7500 535.4350 ;
      RECT 677.4500 532.4350 682.6000 535.4350 ;
      RECT 669.3000 532.4350 674.4500 535.4350 ;
      RECT 661.1500 532.4350 666.3000 535.4350 ;
      RECT 653.0000 532.4350 658.1500 535.4350 ;
      RECT 644.8500 532.4350 650.0000 535.4350 ;
      RECT 636.7000 532.4350 641.8500 535.4350 ;
      RECT 628.5500 532.4350 633.7000 535.4350 ;
      RECT 620.4000 532.4350 625.5500 535.4350 ;
      RECT 612.2500 532.4350 617.4000 535.4350 ;
      RECT 604.1000 532.4350 609.2500 535.4350 ;
      RECT 595.9500 532.4350 601.1000 535.4350 ;
      RECT 587.8000 532.4350 592.9500 535.4350 ;
      RECT 579.6500 532.4350 584.8000 535.4350 ;
      RECT 571.5000 532.4350 576.6500 535.4350 ;
      RECT 563.3500 532.4350 568.5000 535.4350 ;
      RECT 555.2000 532.4350 560.3500 535.4350 ;
      RECT 547.0500 532.4350 552.2000 535.4350 ;
      RECT 538.9000 532.4350 544.0500 535.4350 ;
      RECT 530.7500 532.4350 535.9000 535.4350 ;
      RECT 522.6000 532.4350 527.7500 535.4350 ;
      RECT 514.4500 532.4350 519.6000 535.4350 ;
      RECT 506.3000 532.4350 511.4500 535.4350 ;
      RECT 498.1500 532.4350 503.3000 535.4350 ;
      RECT 490.0000 532.4350 495.1500 535.4350 ;
      RECT 481.8500 532.4350 487.0000 535.4350 ;
      RECT 473.7000 532.4350 478.8500 535.4350 ;
      RECT 465.5500 532.4350 470.7000 535.4350 ;
      RECT 457.4000 532.4350 462.5500 535.4350 ;
      RECT 449.2500 532.4350 454.4000 535.4350 ;
      RECT 441.1000 532.4350 446.2500 535.4350 ;
      RECT 432.9500 532.4350 438.1000 535.4350 ;
      RECT 424.8000 532.4350 429.9500 535.4350 ;
      RECT 416.6500 532.4350 421.8000 535.4350 ;
      RECT 396.5000 532.4350 413.6500 535.4350 ;
      RECT 346.5000 532.4350 393.5000 535.4350 ;
      RECT 326.4650 532.4350 343.5000 535.4350 ;
      RECT 317.9500 532.4350 323.4650 535.4350 ;
      RECT 309.4350 532.4350 314.9500 535.4350 ;
      RECT 300.9200 532.4350 306.4350 535.4350 ;
      RECT 292.4050 532.4350 297.9200 535.4350 ;
      RECT 283.8900 532.4350 289.4050 535.4350 ;
      RECT 275.3750 532.4350 280.8900 535.4350 ;
      RECT 266.8600 532.4350 272.3750 535.4350 ;
      RECT 258.3450 532.4350 263.8600 535.4350 ;
      RECT 249.8300 532.4350 255.3450 535.4350 ;
      RECT 241.3150 532.4350 246.8300 535.4350 ;
      RECT 232.8000 532.4350 238.3150 535.4350 ;
      RECT 224.2850 532.4350 229.8000 535.4350 ;
      RECT 215.7700 532.4350 221.2850 535.4350 ;
      RECT 207.2550 532.4350 212.7700 535.4350 ;
      RECT 198.7400 532.4350 204.2550 535.4350 ;
      RECT 190.2250 532.4350 195.7400 535.4350 ;
      RECT 181.7100 532.4350 187.2250 535.4350 ;
      RECT 173.1950 532.4350 178.7100 535.4350 ;
      RECT 164.6800 532.4350 170.1950 535.4350 ;
      RECT 156.1650 532.4350 161.6800 535.4350 ;
      RECT 147.6500 532.4350 153.1650 535.4350 ;
      RECT 139.1350 532.4350 144.6500 535.4350 ;
      RECT 130.6200 532.4350 136.1350 535.4350 ;
      RECT 122.1050 532.4350 127.6200 535.4350 ;
      RECT 113.5900 532.4350 119.1050 535.4350 ;
      RECT 105.0750 532.4350 110.5900 535.4350 ;
      RECT 96.5600 532.4350 102.0750 535.4350 ;
      RECT 88.0450 532.4350 93.5600 535.4350 ;
      RECT 79.5300 532.4350 85.0450 535.4350 ;
      RECT 71.0150 532.4350 76.5300 535.4350 ;
      RECT 62.5000 532.4350 68.0150 535.4350 ;
      RECT 46.5000 532.4350 59.5000 535.4350 ;
      RECT 8.5000 532.4350 43.5000 535.4350 ;
      RECT 0.0000 532.4350 5.5000 535.4350 ;
      RECT 0.0000 530.9000 1120.0000 532.4350 ;
      RECT 1116.6000 530.4350 1120.0000 530.9000 ;
      RECT 0.0000 528.3400 1113.6000 530.9000 ;
      RECT 1118.5000 527.4350 1120.0000 530.4350 ;
      RECT 1114.5000 525.3400 1120.0000 527.4350 ;
      RECT 1076.5000 525.3400 1111.5000 528.3400 ;
      RECT 1060.5000 525.3400 1073.5000 528.3400 ;
      RECT 1052.3500 525.3400 1057.5000 528.3400 ;
      RECT 1044.2000 525.3400 1049.3500 528.3400 ;
      RECT 1036.0500 525.3400 1041.2000 528.3400 ;
      RECT 1027.9000 525.3400 1033.0500 528.3400 ;
      RECT 1019.7500 525.3400 1024.9000 528.3400 ;
      RECT 1011.6000 525.3400 1016.7500 528.3400 ;
      RECT 1003.4500 525.3400 1008.6000 528.3400 ;
      RECT 995.3000 525.3400 1000.4500 528.3400 ;
      RECT 987.1500 525.3400 992.3000 528.3400 ;
      RECT 979.0000 525.3400 984.1500 528.3400 ;
      RECT 970.8500 525.3400 976.0000 528.3400 ;
      RECT 962.7000 525.3400 967.8500 528.3400 ;
      RECT 954.5500 525.3400 959.7000 528.3400 ;
      RECT 946.4000 525.3400 951.5500 528.3400 ;
      RECT 938.2500 525.3400 943.4000 528.3400 ;
      RECT 930.1000 525.3400 935.2500 528.3400 ;
      RECT 921.9500 525.3400 927.1000 528.3400 ;
      RECT 913.8000 525.3400 918.9500 528.3400 ;
      RECT 905.6500 525.3400 910.8000 528.3400 ;
      RECT 897.5000 525.3400 902.6500 528.3400 ;
      RECT 889.3500 525.3400 894.5000 528.3400 ;
      RECT 881.2000 525.3400 886.3500 528.3400 ;
      RECT 873.0500 525.3400 878.2000 528.3400 ;
      RECT 864.9000 525.3400 870.0500 528.3400 ;
      RECT 856.7500 525.3400 861.9000 528.3400 ;
      RECT 848.6000 525.3400 853.7500 528.3400 ;
      RECT 840.4500 525.3400 845.6000 528.3400 ;
      RECT 832.3000 525.3400 837.4500 528.3400 ;
      RECT 824.1500 525.3400 829.3000 528.3400 ;
      RECT 816.0000 525.3400 821.1500 528.3400 ;
      RECT 807.8500 525.3400 813.0000 528.3400 ;
      RECT 799.7000 525.3400 804.8500 528.3400 ;
      RECT 791.5500 525.3400 796.7000 528.3400 ;
      RECT 783.4000 525.3400 788.5500 528.3400 ;
      RECT 775.2500 525.3400 780.4000 528.3400 ;
      RECT 767.1000 525.3400 772.2500 528.3400 ;
      RECT 758.9500 525.3400 764.1000 528.3400 ;
      RECT 750.8000 525.3400 755.9500 528.3400 ;
      RECT 742.6500 525.3400 747.8000 528.3400 ;
      RECT 734.5000 525.3400 739.6500 528.3400 ;
      RECT 726.3500 525.3400 731.5000 528.3400 ;
      RECT 718.2000 525.3400 723.3500 528.3400 ;
      RECT 710.0500 525.3400 715.2000 528.3400 ;
      RECT 701.9000 525.3400 707.0500 528.3400 ;
      RECT 693.7500 525.3400 698.9000 528.3400 ;
      RECT 685.6000 525.3400 690.7500 528.3400 ;
      RECT 677.4500 525.3400 682.6000 528.3400 ;
      RECT 669.3000 525.3400 674.4500 528.3400 ;
      RECT 661.1500 525.3400 666.3000 528.3400 ;
      RECT 653.0000 525.3400 658.1500 528.3400 ;
      RECT 644.8500 525.3400 650.0000 528.3400 ;
      RECT 636.7000 525.3400 641.8500 528.3400 ;
      RECT 628.5500 525.3400 633.7000 528.3400 ;
      RECT 620.4000 525.3400 625.5500 528.3400 ;
      RECT 612.2500 525.3400 617.4000 528.3400 ;
      RECT 604.1000 525.3400 609.2500 528.3400 ;
      RECT 595.9500 525.3400 601.1000 528.3400 ;
      RECT 587.8000 525.3400 592.9500 528.3400 ;
      RECT 579.6500 525.3400 584.8000 528.3400 ;
      RECT 571.5000 525.3400 576.6500 528.3400 ;
      RECT 563.3500 525.3400 568.5000 528.3400 ;
      RECT 555.2000 525.3400 560.3500 528.3400 ;
      RECT 547.0500 525.3400 552.2000 528.3400 ;
      RECT 538.9000 525.3400 544.0500 528.3400 ;
      RECT 530.7500 525.3400 535.9000 528.3400 ;
      RECT 522.6000 525.3400 527.7500 528.3400 ;
      RECT 514.4500 525.3400 519.6000 528.3400 ;
      RECT 506.3000 525.3400 511.4500 528.3400 ;
      RECT 498.1500 525.3400 503.3000 528.3400 ;
      RECT 490.0000 525.3400 495.1500 528.3400 ;
      RECT 481.8500 525.3400 487.0000 528.3400 ;
      RECT 473.7000 525.3400 478.8500 528.3400 ;
      RECT 465.5500 525.3400 470.7000 528.3400 ;
      RECT 457.4000 525.3400 462.5500 528.3400 ;
      RECT 449.2500 525.3400 454.4000 528.3400 ;
      RECT 441.1000 525.3400 446.2500 528.3400 ;
      RECT 432.9500 525.3400 438.1000 528.3400 ;
      RECT 424.8000 525.3400 429.9500 528.3400 ;
      RECT 416.6500 525.3400 421.8000 528.3400 ;
      RECT 396.5000 525.3400 413.6500 528.3400 ;
      RECT 346.5000 525.3400 393.5000 528.3400 ;
      RECT 326.4650 525.3400 343.5000 528.3400 ;
      RECT 317.9500 525.3400 323.4650 528.3400 ;
      RECT 309.4350 525.3400 314.9500 528.3400 ;
      RECT 300.9200 525.3400 306.4350 528.3400 ;
      RECT 292.4050 525.3400 297.9200 528.3400 ;
      RECT 283.8900 525.3400 289.4050 528.3400 ;
      RECT 275.3750 525.3400 280.8900 528.3400 ;
      RECT 266.8600 525.3400 272.3750 528.3400 ;
      RECT 258.3450 525.3400 263.8600 528.3400 ;
      RECT 249.8300 525.3400 255.3450 528.3400 ;
      RECT 241.3150 525.3400 246.8300 528.3400 ;
      RECT 232.8000 525.3400 238.3150 528.3400 ;
      RECT 224.2850 525.3400 229.8000 528.3400 ;
      RECT 215.7700 525.3400 221.2850 528.3400 ;
      RECT 207.2550 525.3400 212.7700 528.3400 ;
      RECT 198.7400 525.3400 204.2550 528.3400 ;
      RECT 190.2250 525.3400 195.7400 528.3400 ;
      RECT 181.7100 525.3400 187.2250 528.3400 ;
      RECT 173.1950 525.3400 178.7100 528.3400 ;
      RECT 164.6800 525.3400 170.1950 528.3400 ;
      RECT 156.1650 525.3400 161.6800 528.3400 ;
      RECT 147.6500 525.3400 153.1650 528.3400 ;
      RECT 139.1350 525.3400 144.6500 528.3400 ;
      RECT 130.6200 525.3400 136.1350 528.3400 ;
      RECT 122.1050 525.3400 127.6200 528.3400 ;
      RECT 113.5900 525.3400 119.1050 528.3400 ;
      RECT 105.0750 525.3400 110.5900 528.3400 ;
      RECT 96.5600 525.3400 102.0750 528.3400 ;
      RECT 88.0450 525.3400 93.5600 528.3400 ;
      RECT 79.5300 525.3400 85.0450 528.3400 ;
      RECT 71.0150 525.3400 76.5300 528.3400 ;
      RECT 62.5000 525.3400 68.0150 528.3400 ;
      RECT 46.5000 525.3400 59.5000 528.3400 ;
      RECT 8.5000 525.3400 43.5000 528.3400 ;
      RECT 0.0000 525.3400 5.5000 528.3400 ;
      RECT 0.0000 524.5000 1120.0000 525.3400 ;
      RECT 1116.6000 523.3400 1120.0000 524.5000 ;
      RECT 0.0000 521.2450 1113.6000 524.5000 ;
      RECT 1118.5000 520.3400 1120.0000 523.3400 ;
      RECT 1114.5000 518.2450 1120.0000 520.3400 ;
      RECT 1076.5000 518.2450 1111.5000 521.2450 ;
      RECT 1060.5000 518.2450 1073.5000 521.2450 ;
      RECT 1052.3500 518.2450 1057.5000 521.2450 ;
      RECT 1044.2000 518.2450 1049.3500 521.2450 ;
      RECT 1036.0500 518.2450 1041.2000 521.2450 ;
      RECT 1027.9000 518.2450 1033.0500 521.2450 ;
      RECT 1019.7500 518.2450 1024.9000 521.2450 ;
      RECT 1011.6000 518.2450 1016.7500 521.2450 ;
      RECT 1003.4500 518.2450 1008.6000 521.2450 ;
      RECT 995.3000 518.2450 1000.4500 521.2450 ;
      RECT 987.1500 518.2450 992.3000 521.2450 ;
      RECT 979.0000 518.2450 984.1500 521.2450 ;
      RECT 970.8500 518.2450 976.0000 521.2450 ;
      RECT 962.7000 518.2450 967.8500 521.2450 ;
      RECT 954.5500 518.2450 959.7000 521.2450 ;
      RECT 946.4000 518.2450 951.5500 521.2450 ;
      RECT 938.2500 518.2450 943.4000 521.2450 ;
      RECT 930.1000 518.2450 935.2500 521.2450 ;
      RECT 921.9500 518.2450 927.1000 521.2450 ;
      RECT 913.8000 518.2450 918.9500 521.2450 ;
      RECT 905.6500 518.2450 910.8000 521.2450 ;
      RECT 897.5000 518.2450 902.6500 521.2450 ;
      RECT 889.3500 518.2450 894.5000 521.2450 ;
      RECT 881.2000 518.2450 886.3500 521.2450 ;
      RECT 873.0500 518.2450 878.2000 521.2450 ;
      RECT 864.9000 518.2450 870.0500 521.2450 ;
      RECT 856.7500 518.2450 861.9000 521.2450 ;
      RECT 848.6000 518.2450 853.7500 521.2450 ;
      RECT 840.4500 518.2450 845.6000 521.2450 ;
      RECT 832.3000 518.2450 837.4500 521.2450 ;
      RECT 824.1500 518.2450 829.3000 521.2450 ;
      RECT 816.0000 518.2450 821.1500 521.2450 ;
      RECT 807.8500 518.2450 813.0000 521.2450 ;
      RECT 799.7000 518.2450 804.8500 521.2450 ;
      RECT 791.5500 518.2450 796.7000 521.2450 ;
      RECT 783.4000 518.2450 788.5500 521.2450 ;
      RECT 775.2500 518.2450 780.4000 521.2450 ;
      RECT 767.1000 518.2450 772.2500 521.2450 ;
      RECT 758.9500 518.2450 764.1000 521.2450 ;
      RECT 750.8000 518.2450 755.9500 521.2450 ;
      RECT 742.6500 518.2450 747.8000 521.2450 ;
      RECT 734.5000 518.2450 739.6500 521.2450 ;
      RECT 726.3500 518.2450 731.5000 521.2450 ;
      RECT 718.2000 518.2450 723.3500 521.2450 ;
      RECT 710.0500 518.2450 715.2000 521.2450 ;
      RECT 701.9000 518.2450 707.0500 521.2450 ;
      RECT 693.7500 518.2450 698.9000 521.2450 ;
      RECT 685.6000 518.2450 690.7500 521.2450 ;
      RECT 677.4500 518.2450 682.6000 521.2450 ;
      RECT 669.3000 518.2450 674.4500 521.2450 ;
      RECT 661.1500 518.2450 666.3000 521.2450 ;
      RECT 653.0000 518.2450 658.1500 521.2450 ;
      RECT 644.8500 518.2450 650.0000 521.2450 ;
      RECT 636.7000 518.2450 641.8500 521.2450 ;
      RECT 628.5500 518.2450 633.7000 521.2450 ;
      RECT 620.4000 518.2450 625.5500 521.2450 ;
      RECT 612.2500 518.2450 617.4000 521.2450 ;
      RECT 604.1000 518.2450 609.2500 521.2450 ;
      RECT 595.9500 518.2450 601.1000 521.2450 ;
      RECT 587.8000 518.2450 592.9500 521.2450 ;
      RECT 579.6500 518.2450 584.8000 521.2450 ;
      RECT 571.5000 518.2450 576.6500 521.2450 ;
      RECT 563.3500 518.2450 568.5000 521.2450 ;
      RECT 555.2000 518.2450 560.3500 521.2450 ;
      RECT 547.0500 518.2450 552.2000 521.2450 ;
      RECT 538.9000 518.2450 544.0500 521.2450 ;
      RECT 530.7500 518.2450 535.9000 521.2450 ;
      RECT 522.6000 518.2450 527.7500 521.2450 ;
      RECT 514.4500 518.2450 519.6000 521.2450 ;
      RECT 506.3000 518.2450 511.4500 521.2450 ;
      RECT 498.1500 518.2450 503.3000 521.2450 ;
      RECT 490.0000 518.2450 495.1500 521.2450 ;
      RECT 481.8500 518.2450 487.0000 521.2450 ;
      RECT 473.7000 518.2450 478.8500 521.2450 ;
      RECT 465.5500 518.2450 470.7000 521.2450 ;
      RECT 457.4000 518.2450 462.5500 521.2450 ;
      RECT 449.2500 518.2450 454.4000 521.2450 ;
      RECT 441.1000 518.2450 446.2500 521.2450 ;
      RECT 432.9500 518.2450 438.1000 521.2450 ;
      RECT 424.8000 518.2450 429.9500 521.2450 ;
      RECT 416.6500 518.2450 421.8000 521.2450 ;
      RECT 396.5000 518.2450 413.6500 521.2450 ;
      RECT 346.5000 518.2450 393.5000 521.2450 ;
      RECT 326.4650 518.2450 343.5000 521.2450 ;
      RECT 317.9500 518.2450 323.4650 521.2450 ;
      RECT 309.4350 518.2450 314.9500 521.2450 ;
      RECT 300.9200 518.2450 306.4350 521.2450 ;
      RECT 292.4050 518.2450 297.9200 521.2450 ;
      RECT 283.8900 518.2450 289.4050 521.2450 ;
      RECT 275.3750 518.2450 280.8900 521.2450 ;
      RECT 266.8600 518.2450 272.3750 521.2450 ;
      RECT 258.3450 518.2450 263.8600 521.2450 ;
      RECT 249.8300 518.2450 255.3450 521.2450 ;
      RECT 241.3150 518.2450 246.8300 521.2450 ;
      RECT 232.8000 518.2450 238.3150 521.2450 ;
      RECT 224.2850 518.2450 229.8000 521.2450 ;
      RECT 215.7700 518.2450 221.2850 521.2450 ;
      RECT 207.2550 518.2450 212.7700 521.2450 ;
      RECT 198.7400 518.2450 204.2550 521.2450 ;
      RECT 190.2250 518.2450 195.7400 521.2450 ;
      RECT 181.7100 518.2450 187.2250 521.2450 ;
      RECT 173.1950 518.2450 178.7100 521.2450 ;
      RECT 164.6800 518.2450 170.1950 521.2450 ;
      RECT 156.1650 518.2450 161.6800 521.2450 ;
      RECT 147.6500 518.2450 153.1650 521.2450 ;
      RECT 139.1350 518.2450 144.6500 521.2450 ;
      RECT 130.6200 518.2450 136.1350 521.2450 ;
      RECT 122.1050 518.2450 127.6200 521.2450 ;
      RECT 113.5900 518.2450 119.1050 521.2450 ;
      RECT 105.0750 518.2450 110.5900 521.2450 ;
      RECT 96.5600 518.2450 102.0750 521.2450 ;
      RECT 88.0450 518.2450 93.5600 521.2450 ;
      RECT 79.5300 518.2450 85.0450 521.2450 ;
      RECT 71.0150 518.2450 76.5300 521.2450 ;
      RECT 62.5000 518.2450 68.0150 521.2450 ;
      RECT 46.5000 518.2450 59.5000 521.2450 ;
      RECT 8.5000 518.2450 43.5000 521.2450 ;
      RECT 0.0000 518.2450 5.5000 521.2450 ;
      RECT 0.0000 517.3000 1120.0000 518.2450 ;
      RECT 1116.6000 516.2450 1120.0000 517.3000 ;
      RECT 0.0000 514.1500 1113.6000 517.3000 ;
      RECT 1118.5000 513.2450 1120.0000 516.2450 ;
      RECT 1114.5000 511.1500 1120.0000 513.2450 ;
      RECT 1076.5000 511.1500 1111.5000 514.1500 ;
      RECT 1060.5000 511.1500 1073.5000 514.1500 ;
      RECT 1052.3500 511.1500 1057.5000 514.1500 ;
      RECT 1044.2000 511.1500 1049.3500 514.1500 ;
      RECT 1036.0500 511.1500 1041.2000 514.1500 ;
      RECT 1027.9000 511.1500 1033.0500 514.1500 ;
      RECT 1019.7500 511.1500 1024.9000 514.1500 ;
      RECT 1011.6000 511.1500 1016.7500 514.1500 ;
      RECT 1003.4500 511.1500 1008.6000 514.1500 ;
      RECT 995.3000 511.1500 1000.4500 514.1500 ;
      RECT 987.1500 511.1500 992.3000 514.1500 ;
      RECT 979.0000 511.1500 984.1500 514.1500 ;
      RECT 970.8500 511.1500 976.0000 514.1500 ;
      RECT 962.7000 511.1500 967.8500 514.1500 ;
      RECT 954.5500 511.1500 959.7000 514.1500 ;
      RECT 946.4000 511.1500 951.5500 514.1500 ;
      RECT 938.2500 511.1500 943.4000 514.1500 ;
      RECT 930.1000 511.1500 935.2500 514.1500 ;
      RECT 921.9500 511.1500 927.1000 514.1500 ;
      RECT 913.8000 511.1500 918.9500 514.1500 ;
      RECT 905.6500 511.1500 910.8000 514.1500 ;
      RECT 897.5000 511.1500 902.6500 514.1500 ;
      RECT 889.3500 511.1500 894.5000 514.1500 ;
      RECT 881.2000 511.1500 886.3500 514.1500 ;
      RECT 873.0500 511.1500 878.2000 514.1500 ;
      RECT 864.9000 511.1500 870.0500 514.1500 ;
      RECT 856.7500 511.1500 861.9000 514.1500 ;
      RECT 848.6000 511.1500 853.7500 514.1500 ;
      RECT 840.4500 511.1500 845.6000 514.1500 ;
      RECT 832.3000 511.1500 837.4500 514.1500 ;
      RECT 824.1500 511.1500 829.3000 514.1500 ;
      RECT 816.0000 511.1500 821.1500 514.1500 ;
      RECT 807.8500 511.1500 813.0000 514.1500 ;
      RECT 799.7000 511.1500 804.8500 514.1500 ;
      RECT 791.5500 511.1500 796.7000 514.1500 ;
      RECT 783.4000 511.1500 788.5500 514.1500 ;
      RECT 775.2500 511.1500 780.4000 514.1500 ;
      RECT 767.1000 511.1500 772.2500 514.1500 ;
      RECT 758.9500 511.1500 764.1000 514.1500 ;
      RECT 750.8000 511.1500 755.9500 514.1500 ;
      RECT 742.6500 511.1500 747.8000 514.1500 ;
      RECT 734.5000 511.1500 739.6500 514.1500 ;
      RECT 726.3500 511.1500 731.5000 514.1500 ;
      RECT 718.2000 511.1500 723.3500 514.1500 ;
      RECT 710.0500 511.1500 715.2000 514.1500 ;
      RECT 701.9000 511.1500 707.0500 514.1500 ;
      RECT 693.7500 511.1500 698.9000 514.1500 ;
      RECT 685.6000 511.1500 690.7500 514.1500 ;
      RECT 677.4500 511.1500 682.6000 514.1500 ;
      RECT 669.3000 511.1500 674.4500 514.1500 ;
      RECT 661.1500 511.1500 666.3000 514.1500 ;
      RECT 653.0000 511.1500 658.1500 514.1500 ;
      RECT 644.8500 511.1500 650.0000 514.1500 ;
      RECT 636.7000 511.1500 641.8500 514.1500 ;
      RECT 628.5500 511.1500 633.7000 514.1500 ;
      RECT 620.4000 511.1500 625.5500 514.1500 ;
      RECT 612.2500 511.1500 617.4000 514.1500 ;
      RECT 604.1000 511.1500 609.2500 514.1500 ;
      RECT 595.9500 511.1500 601.1000 514.1500 ;
      RECT 587.8000 511.1500 592.9500 514.1500 ;
      RECT 579.6500 511.1500 584.8000 514.1500 ;
      RECT 571.5000 511.1500 576.6500 514.1500 ;
      RECT 563.3500 511.1500 568.5000 514.1500 ;
      RECT 555.2000 511.1500 560.3500 514.1500 ;
      RECT 547.0500 511.1500 552.2000 514.1500 ;
      RECT 538.9000 511.1500 544.0500 514.1500 ;
      RECT 530.7500 511.1500 535.9000 514.1500 ;
      RECT 522.6000 511.1500 527.7500 514.1500 ;
      RECT 514.4500 511.1500 519.6000 514.1500 ;
      RECT 506.3000 511.1500 511.4500 514.1500 ;
      RECT 498.1500 511.1500 503.3000 514.1500 ;
      RECT 490.0000 511.1500 495.1500 514.1500 ;
      RECT 481.8500 511.1500 487.0000 514.1500 ;
      RECT 473.7000 511.1500 478.8500 514.1500 ;
      RECT 465.5500 511.1500 470.7000 514.1500 ;
      RECT 457.4000 511.1500 462.5500 514.1500 ;
      RECT 449.2500 511.1500 454.4000 514.1500 ;
      RECT 441.1000 511.1500 446.2500 514.1500 ;
      RECT 432.9500 511.1500 438.1000 514.1500 ;
      RECT 424.8000 511.1500 429.9500 514.1500 ;
      RECT 416.6500 511.1500 421.8000 514.1500 ;
      RECT 396.5000 511.1500 413.6500 514.1500 ;
      RECT 346.5000 511.1500 393.5000 514.1500 ;
      RECT 326.4650 511.1500 343.5000 514.1500 ;
      RECT 317.9500 511.1500 323.4650 514.1500 ;
      RECT 309.4350 511.1500 314.9500 514.1500 ;
      RECT 300.9200 511.1500 306.4350 514.1500 ;
      RECT 292.4050 511.1500 297.9200 514.1500 ;
      RECT 283.8900 511.1500 289.4050 514.1500 ;
      RECT 275.3750 511.1500 280.8900 514.1500 ;
      RECT 266.8600 511.1500 272.3750 514.1500 ;
      RECT 258.3450 511.1500 263.8600 514.1500 ;
      RECT 249.8300 511.1500 255.3450 514.1500 ;
      RECT 241.3150 511.1500 246.8300 514.1500 ;
      RECT 232.8000 511.1500 238.3150 514.1500 ;
      RECT 224.2850 511.1500 229.8000 514.1500 ;
      RECT 215.7700 511.1500 221.2850 514.1500 ;
      RECT 207.2550 511.1500 212.7700 514.1500 ;
      RECT 198.7400 511.1500 204.2550 514.1500 ;
      RECT 190.2250 511.1500 195.7400 514.1500 ;
      RECT 181.7100 511.1500 187.2250 514.1500 ;
      RECT 173.1950 511.1500 178.7100 514.1500 ;
      RECT 164.6800 511.1500 170.1950 514.1500 ;
      RECT 156.1650 511.1500 161.6800 514.1500 ;
      RECT 147.6500 511.1500 153.1650 514.1500 ;
      RECT 139.1350 511.1500 144.6500 514.1500 ;
      RECT 130.6200 511.1500 136.1350 514.1500 ;
      RECT 122.1050 511.1500 127.6200 514.1500 ;
      RECT 113.5900 511.1500 119.1050 514.1500 ;
      RECT 105.0750 511.1500 110.5900 514.1500 ;
      RECT 96.5600 511.1500 102.0750 514.1500 ;
      RECT 88.0450 511.1500 93.5600 514.1500 ;
      RECT 79.5300 511.1500 85.0450 514.1500 ;
      RECT 71.0150 511.1500 76.5300 514.1500 ;
      RECT 62.5000 511.1500 68.0150 514.1500 ;
      RECT 46.5000 511.1500 59.5000 514.1500 ;
      RECT 8.5000 511.1500 43.5000 514.1500 ;
      RECT 0.0000 511.1500 5.5000 514.1500 ;
      RECT 0.0000 509.7000 1120.0000 511.1500 ;
      RECT 1116.6000 509.1500 1120.0000 509.7000 ;
      RECT 0.0000 507.0550 1113.6000 509.7000 ;
      RECT 1118.5000 506.1500 1120.0000 509.1500 ;
      RECT 1114.5000 504.0550 1120.0000 506.1500 ;
      RECT 1076.5000 504.0550 1111.5000 507.0550 ;
      RECT 1060.5000 504.0550 1073.5000 507.0550 ;
      RECT 1052.3500 504.0550 1057.5000 507.0550 ;
      RECT 1044.2000 504.0550 1049.3500 507.0550 ;
      RECT 1036.0500 504.0550 1041.2000 507.0550 ;
      RECT 1027.9000 504.0550 1033.0500 507.0550 ;
      RECT 1019.7500 504.0550 1024.9000 507.0550 ;
      RECT 1011.6000 504.0550 1016.7500 507.0550 ;
      RECT 1003.4500 504.0550 1008.6000 507.0550 ;
      RECT 995.3000 504.0550 1000.4500 507.0550 ;
      RECT 987.1500 504.0550 992.3000 507.0550 ;
      RECT 979.0000 504.0550 984.1500 507.0550 ;
      RECT 970.8500 504.0550 976.0000 507.0550 ;
      RECT 962.7000 504.0550 967.8500 507.0550 ;
      RECT 954.5500 504.0550 959.7000 507.0550 ;
      RECT 946.4000 504.0550 951.5500 507.0550 ;
      RECT 938.2500 504.0550 943.4000 507.0550 ;
      RECT 930.1000 504.0550 935.2500 507.0550 ;
      RECT 921.9500 504.0550 927.1000 507.0550 ;
      RECT 913.8000 504.0550 918.9500 507.0550 ;
      RECT 905.6500 504.0550 910.8000 507.0550 ;
      RECT 897.5000 504.0550 902.6500 507.0550 ;
      RECT 889.3500 504.0550 894.5000 507.0550 ;
      RECT 881.2000 504.0550 886.3500 507.0550 ;
      RECT 873.0500 504.0550 878.2000 507.0550 ;
      RECT 864.9000 504.0550 870.0500 507.0550 ;
      RECT 856.7500 504.0550 861.9000 507.0550 ;
      RECT 848.6000 504.0550 853.7500 507.0550 ;
      RECT 840.4500 504.0550 845.6000 507.0550 ;
      RECT 832.3000 504.0550 837.4500 507.0550 ;
      RECT 824.1500 504.0550 829.3000 507.0550 ;
      RECT 816.0000 504.0550 821.1500 507.0550 ;
      RECT 807.8500 504.0550 813.0000 507.0550 ;
      RECT 799.7000 504.0550 804.8500 507.0550 ;
      RECT 791.5500 504.0550 796.7000 507.0550 ;
      RECT 783.4000 504.0550 788.5500 507.0550 ;
      RECT 775.2500 504.0550 780.4000 507.0550 ;
      RECT 767.1000 504.0550 772.2500 507.0550 ;
      RECT 758.9500 504.0550 764.1000 507.0550 ;
      RECT 750.8000 504.0550 755.9500 507.0550 ;
      RECT 742.6500 504.0550 747.8000 507.0550 ;
      RECT 734.5000 504.0550 739.6500 507.0550 ;
      RECT 726.3500 504.0550 731.5000 507.0550 ;
      RECT 718.2000 504.0550 723.3500 507.0550 ;
      RECT 710.0500 504.0550 715.2000 507.0550 ;
      RECT 701.9000 504.0550 707.0500 507.0550 ;
      RECT 693.7500 504.0550 698.9000 507.0550 ;
      RECT 685.6000 504.0550 690.7500 507.0550 ;
      RECT 677.4500 504.0550 682.6000 507.0550 ;
      RECT 669.3000 504.0550 674.4500 507.0550 ;
      RECT 661.1500 504.0550 666.3000 507.0550 ;
      RECT 653.0000 504.0550 658.1500 507.0550 ;
      RECT 644.8500 504.0550 650.0000 507.0550 ;
      RECT 636.7000 504.0550 641.8500 507.0550 ;
      RECT 628.5500 504.0550 633.7000 507.0550 ;
      RECT 620.4000 504.0550 625.5500 507.0550 ;
      RECT 612.2500 504.0550 617.4000 507.0550 ;
      RECT 604.1000 504.0550 609.2500 507.0550 ;
      RECT 595.9500 504.0550 601.1000 507.0550 ;
      RECT 587.8000 504.0550 592.9500 507.0550 ;
      RECT 579.6500 504.0550 584.8000 507.0550 ;
      RECT 571.5000 504.0550 576.6500 507.0550 ;
      RECT 563.3500 504.0550 568.5000 507.0550 ;
      RECT 555.2000 504.0550 560.3500 507.0550 ;
      RECT 547.0500 504.0550 552.2000 507.0550 ;
      RECT 538.9000 504.0550 544.0500 507.0550 ;
      RECT 530.7500 504.0550 535.9000 507.0550 ;
      RECT 522.6000 504.0550 527.7500 507.0550 ;
      RECT 514.4500 504.0550 519.6000 507.0550 ;
      RECT 506.3000 504.0550 511.4500 507.0550 ;
      RECT 498.1500 504.0550 503.3000 507.0550 ;
      RECT 490.0000 504.0550 495.1500 507.0550 ;
      RECT 481.8500 504.0550 487.0000 507.0550 ;
      RECT 473.7000 504.0550 478.8500 507.0550 ;
      RECT 465.5500 504.0550 470.7000 507.0550 ;
      RECT 457.4000 504.0550 462.5500 507.0550 ;
      RECT 449.2500 504.0550 454.4000 507.0550 ;
      RECT 441.1000 504.0550 446.2500 507.0550 ;
      RECT 432.9500 504.0550 438.1000 507.0550 ;
      RECT 424.8000 504.0550 429.9500 507.0550 ;
      RECT 416.6500 504.0550 421.8000 507.0550 ;
      RECT 396.5000 504.0550 413.6500 507.0550 ;
      RECT 346.5000 504.0550 393.5000 507.0550 ;
      RECT 326.4650 504.0550 343.5000 507.0550 ;
      RECT 317.9500 504.0550 323.4650 507.0550 ;
      RECT 309.4350 504.0550 314.9500 507.0550 ;
      RECT 300.9200 504.0550 306.4350 507.0550 ;
      RECT 292.4050 504.0550 297.9200 507.0550 ;
      RECT 283.8900 504.0550 289.4050 507.0550 ;
      RECT 275.3750 504.0550 280.8900 507.0550 ;
      RECT 266.8600 504.0550 272.3750 507.0550 ;
      RECT 258.3450 504.0550 263.8600 507.0550 ;
      RECT 249.8300 504.0550 255.3450 507.0550 ;
      RECT 241.3150 504.0550 246.8300 507.0550 ;
      RECT 232.8000 504.0550 238.3150 507.0550 ;
      RECT 224.2850 504.0550 229.8000 507.0550 ;
      RECT 215.7700 504.0550 221.2850 507.0550 ;
      RECT 207.2550 504.0550 212.7700 507.0550 ;
      RECT 198.7400 504.0550 204.2550 507.0550 ;
      RECT 190.2250 504.0550 195.7400 507.0550 ;
      RECT 181.7100 504.0550 187.2250 507.0550 ;
      RECT 173.1950 504.0550 178.7100 507.0550 ;
      RECT 164.6800 504.0550 170.1950 507.0550 ;
      RECT 156.1650 504.0550 161.6800 507.0550 ;
      RECT 147.6500 504.0550 153.1650 507.0550 ;
      RECT 139.1350 504.0550 144.6500 507.0550 ;
      RECT 130.6200 504.0550 136.1350 507.0550 ;
      RECT 122.1050 504.0550 127.6200 507.0550 ;
      RECT 113.5900 504.0550 119.1050 507.0550 ;
      RECT 105.0750 504.0550 110.5900 507.0550 ;
      RECT 96.5600 504.0550 102.0750 507.0550 ;
      RECT 88.0450 504.0550 93.5600 507.0550 ;
      RECT 79.5300 504.0550 85.0450 507.0550 ;
      RECT 71.0150 504.0550 76.5300 507.0550 ;
      RECT 62.5000 504.0550 68.0150 507.0550 ;
      RECT 46.5000 504.0550 59.5000 507.0550 ;
      RECT 8.5000 504.0550 43.5000 507.0550 ;
      RECT 0.0000 504.0550 5.5000 507.0550 ;
      RECT 0.0000 502.5000 1120.0000 504.0550 ;
      RECT 1116.6000 502.0550 1120.0000 502.5000 ;
      RECT 0.0000 499.9600 1113.6000 502.5000 ;
      RECT 1118.5000 499.0550 1120.0000 502.0550 ;
      RECT 1114.5000 496.9600 1120.0000 499.0550 ;
      RECT 1076.5000 496.9600 1111.5000 499.9600 ;
      RECT 1060.5000 496.9600 1073.5000 499.9600 ;
      RECT 1052.3500 496.9600 1057.5000 499.9600 ;
      RECT 1044.2000 496.9600 1049.3500 499.9600 ;
      RECT 1036.0500 496.9600 1041.2000 499.9600 ;
      RECT 1027.9000 496.9600 1033.0500 499.9600 ;
      RECT 1019.7500 496.9600 1024.9000 499.9600 ;
      RECT 1011.6000 496.9600 1016.7500 499.9600 ;
      RECT 1003.4500 496.9600 1008.6000 499.9600 ;
      RECT 995.3000 496.9600 1000.4500 499.9600 ;
      RECT 987.1500 496.9600 992.3000 499.9600 ;
      RECT 979.0000 496.9600 984.1500 499.9600 ;
      RECT 970.8500 496.9600 976.0000 499.9600 ;
      RECT 962.7000 496.9600 967.8500 499.9600 ;
      RECT 954.5500 496.9600 959.7000 499.9600 ;
      RECT 946.4000 496.9600 951.5500 499.9600 ;
      RECT 938.2500 496.9600 943.4000 499.9600 ;
      RECT 930.1000 496.9600 935.2500 499.9600 ;
      RECT 921.9500 496.9600 927.1000 499.9600 ;
      RECT 913.8000 496.9600 918.9500 499.9600 ;
      RECT 905.6500 496.9600 910.8000 499.9600 ;
      RECT 897.5000 496.9600 902.6500 499.9600 ;
      RECT 889.3500 496.9600 894.5000 499.9600 ;
      RECT 881.2000 496.9600 886.3500 499.9600 ;
      RECT 873.0500 496.9600 878.2000 499.9600 ;
      RECT 864.9000 496.9600 870.0500 499.9600 ;
      RECT 856.7500 496.9600 861.9000 499.9600 ;
      RECT 848.6000 496.9600 853.7500 499.9600 ;
      RECT 840.4500 496.9600 845.6000 499.9600 ;
      RECT 832.3000 496.9600 837.4500 499.9600 ;
      RECT 824.1500 496.9600 829.3000 499.9600 ;
      RECT 816.0000 496.9600 821.1500 499.9600 ;
      RECT 807.8500 496.9600 813.0000 499.9600 ;
      RECT 799.7000 496.9600 804.8500 499.9600 ;
      RECT 791.5500 496.9600 796.7000 499.9600 ;
      RECT 783.4000 496.9600 788.5500 499.9600 ;
      RECT 775.2500 496.9600 780.4000 499.9600 ;
      RECT 767.1000 496.9600 772.2500 499.9600 ;
      RECT 758.9500 496.9600 764.1000 499.9600 ;
      RECT 750.8000 496.9600 755.9500 499.9600 ;
      RECT 742.6500 496.9600 747.8000 499.9600 ;
      RECT 734.5000 496.9600 739.6500 499.9600 ;
      RECT 726.3500 496.9600 731.5000 499.9600 ;
      RECT 718.2000 496.9600 723.3500 499.9600 ;
      RECT 710.0500 496.9600 715.2000 499.9600 ;
      RECT 701.9000 496.9600 707.0500 499.9600 ;
      RECT 693.7500 496.9600 698.9000 499.9600 ;
      RECT 685.6000 496.9600 690.7500 499.9600 ;
      RECT 677.4500 496.9600 682.6000 499.9600 ;
      RECT 669.3000 496.9600 674.4500 499.9600 ;
      RECT 661.1500 496.9600 666.3000 499.9600 ;
      RECT 653.0000 496.9600 658.1500 499.9600 ;
      RECT 644.8500 496.9600 650.0000 499.9600 ;
      RECT 636.7000 496.9600 641.8500 499.9600 ;
      RECT 628.5500 496.9600 633.7000 499.9600 ;
      RECT 620.4000 496.9600 625.5500 499.9600 ;
      RECT 612.2500 496.9600 617.4000 499.9600 ;
      RECT 604.1000 496.9600 609.2500 499.9600 ;
      RECT 595.9500 496.9600 601.1000 499.9600 ;
      RECT 587.8000 496.9600 592.9500 499.9600 ;
      RECT 579.6500 496.9600 584.8000 499.9600 ;
      RECT 571.5000 496.9600 576.6500 499.9600 ;
      RECT 563.3500 496.9600 568.5000 499.9600 ;
      RECT 555.2000 496.9600 560.3500 499.9600 ;
      RECT 547.0500 496.9600 552.2000 499.9600 ;
      RECT 538.9000 496.9600 544.0500 499.9600 ;
      RECT 530.7500 496.9600 535.9000 499.9600 ;
      RECT 522.6000 496.9600 527.7500 499.9600 ;
      RECT 514.4500 496.9600 519.6000 499.9600 ;
      RECT 506.3000 496.9600 511.4500 499.9600 ;
      RECT 498.1500 496.9600 503.3000 499.9600 ;
      RECT 490.0000 496.9600 495.1500 499.9600 ;
      RECT 481.8500 496.9600 487.0000 499.9600 ;
      RECT 473.7000 496.9600 478.8500 499.9600 ;
      RECT 465.5500 496.9600 470.7000 499.9600 ;
      RECT 457.4000 496.9600 462.5500 499.9600 ;
      RECT 449.2500 496.9600 454.4000 499.9600 ;
      RECT 441.1000 496.9600 446.2500 499.9600 ;
      RECT 432.9500 496.9600 438.1000 499.9600 ;
      RECT 424.8000 496.9600 429.9500 499.9600 ;
      RECT 416.6500 496.9600 421.8000 499.9600 ;
      RECT 396.5000 496.9600 413.6500 499.9600 ;
      RECT 346.5000 496.9600 393.5000 499.9600 ;
      RECT 326.4650 496.9600 343.5000 499.9600 ;
      RECT 317.9500 496.9600 323.4650 499.9600 ;
      RECT 309.4350 496.9600 314.9500 499.9600 ;
      RECT 300.9200 496.9600 306.4350 499.9600 ;
      RECT 292.4050 496.9600 297.9200 499.9600 ;
      RECT 283.8900 496.9600 289.4050 499.9600 ;
      RECT 275.3750 496.9600 280.8900 499.9600 ;
      RECT 266.8600 496.9600 272.3750 499.9600 ;
      RECT 258.3450 496.9600 263.8600 499.9600 ;
      RECT 249.8300 496.9600 255.3450 499.9600 ;
      RECT 241.3150 496.9600 246.8300 499.9600 ;
      RECT 232.8000 496.9600 238.3150 499.9600 ;
      RECT 224.2850 496.9600 229.8000 499.9600 ;
      RECT 215.7700 496.9600 221.2850 499.9600 ;
      RECT 207.2550 496.9600 212.7700 499.9600 ;
      RECT 198.7400 496.9600 204.2550 499.9600 ;
      RECT 190.2250 496.9600 195.7400 499.9600 ;
      RECT 181.7100 496.9600 187.2250 499.9600 ;
      RECT 173.1950 496.9600 178.7100 499.9600 ;
      RECT 164.6800 496.9600 170.1950 499.9600 ;
      RECT 156.1650 496.9600 161.6800 499.9600 ;
      RECT 147.6500 496.9600 153.1650 499.9600 ;
      RECT 139.1350 496.9600 144.6500 499.9600 ;
      RECT 130.6200 496.9600 136.1350 499.9600 ;
      RECT 122.1050 496.9600 127.6200 499.9600 ;
      RECT 113.5900 496.9600 119.1050 499.9600 ;
      RECT 105.0750 496.9600 110.5900 499.9600 ;
      RECT 96.5600 496.9600 102.0750 499.9600 ;
      RECT 88.0450 496.9600 93.5600 499.9600 ;
      RECT 79.5300 496.9600 85.0450 499.9600 ;
      RECT 71.0150 496.9600 76.5300 499.9600 ;
      RECT 62.5000 496.9600 68.0150 499.9600 ;
      RECT 46.5000 496.9600 59.5000 499.9600 ;
      RECT 8.5000 496.9600 43.5000 499.9600 ;
      RECT 0.0000 496.9600 5.5000 499.9600 ;
      RECT 0.0000 495.5000 1120.0000 496.9600 ;
      RECT 1116.6000 494.9600 1120.0000 495.5000 ;
      RECT 0.0000 492.8650 1113.6000 495.5000 ;
      RECT 1118.5000 491.9600 1120.0000 494.9600 ;
      RECT 1114.5000 489.8650 1120.0000 491.9600 ;
      RECT 1076.5000 489.8650 1111.5000 492.8650 ;
      RECT 1060.5000 489.8650 1073.5000 492.8650 ;
      RECT 1052.3500 489.8650 1057.5000 492.8650 ;
      RECT 1044.2000 489.8650 1049.3500 492.8650 ;
      RECT 1036.0500 489.8650 1041.2000 492.8650 ;
      RECT 1027.9000 489.8650 1033.0500 492.8650 ;
      RECT 1019.7500 489.8650 1024.9000 492.8650 ;
      RECT 1011.6000 489.8650 1016.7500 492.8650 ;
      RECT 1003.4500 489.8650 1008.6000 492.8650 ;
      RECT 995.3000 489.8650 1000.4500 492.8650 ;
      RECT 987.1500 489.8650 992.3000 492.8650 ;
      RECT 979.0000 489.8650 984.1500 492.8650 ;
      RECT 970.8500 489.8650 976.0000 492.8650 ;
      RECT 962.7000 489.8650 967.8500 492.8650 ;
      RECT 954.5500 489.8650 959.7000 492.8650 ;
      RECT 946.4000 489.8650 951.5500 492.8650 ;
      RECT 938.2500 489.8650 943.4000 492.8650 ;
      RECT 930.1000 489.8650 935.2500 492.8650 ;
      RECT 921.9500 489.8650 927.1000 492.8650 ;
      RECT 913.8000 489.8650 918.9500 492.8650 ;
      RECT 905.6500 489.8650 910.8000 492.8650 ;
      RECT 897.5000 489.8650 902.6500 492.8650 ;
      RECT 889.3500 489.8650 894.5000 492.8650 ;
      RECT 881.2000 489.8650 886.3500 492.8650 ;
      RECT 873.0500 489.8650 878.2000 492.8650 ;
      RECT 864.9000 489.8650 870.0500 492.8650 ;
      RECT 856.7500 489.8650 861.9000 492.8650 ;
      RECT 848.6000 489.8650 853.7500 492.8650 ;
      RECT 840.4500 489.8650 845.6000 492.8650 ;
      RECT 832.3000 489.8650 837.4500 492.8650 ;
      RECT 824.1500 489.8650 829.3000 492.8650 ;
      RECT 816.0000 489.8650 821.1500 492.8650 ;
      RECT 807.8500 489.8650 813.0000 492.8650 ;
      RECT 799.7000 489.8650 804.8500 492.8650 ;
      RECT 791.5500 489.8650 796.7000 492.8650 ;
      RECT 783.4000 489.8650 788.5500 492.8650 ;
      RECT 775.2500 489.8650 780.4000 492.8650 ;
      RECT 767.1000 489.8650 772.2500 492.8650 ;
      RECT 758.9500 489.8650 764.1000 492.8650 ;
      RECT 750.8000 489.8650 755.9500 492.8650 ;
      RECT 742.6500 489.8650 747.8000 492.8650 ;
      RECT 734.5000 489.8650 739.6500 492.8650 ;
      RECT 726.3500 489.8650 731.5000 492.8650 ;
      RECT 718.2000 489.8650 723.3500 492.8650 ;
      RECT 710.0500 489.8650 715.2000 492.8650 ;
      RECT 701.9000 489.8650 707.0500 492.8650 ;
      RECT 693.7500 489.8650 698.9000 492.8650 ;
      RECT 685.6000 489.8650 690.7500 492.8650 ;
      RECT 677.4500 489.8650 682.6000 492.8650 ;
      RECT 669.3000 489.8650 674.4500 492.8650 ;
      RECT 661.1500 489.8650 666.3000 492.8650 ;
      RECT 653.0000 489.8650 658.1500 492.8650 ;
      RECT 644.8500 489.8650 650.0000 492.8650 ;
      RECT 636.7000 489.8650 641.8500 492.8650 ;
      RECT 628.5500 489.8650 633.7000 492.8650 ;
      RECT 620.4000 489.8650 625.5500 492.8650 ;
      RECT 612.2500 489.8650 617.4000 492.8650 ;
      RECT 604.1000 489.8650 609.2500 492.8650 ;
      RECT 595.9500 489.8650 601.1000 492.8650 ;
      RECT 587.8000 489.8650 592.9500 492.8650 ;
      RECT 579.6500 489.8650 584.8000 492.8650 ;
      RECT 571.5000 489.8650 576.6500 492.8650 ;
      RECT 563.3500 489.8650 568.5000 492.8650 ;
      RECT 555.2000 489.8650 560.3500 492.8650 ;
      RECT 547.0500 489.8650 552.2000 492.8650 ;
      RECT 538.9000 489.8650 544.0500 492.8650 ;
      RECT 530.7500 489.8650 535.9000 492.8650 ;
      RECT 522.6000 489.8650 527.7500 492.8650 ;
      RECT 514.4500 489.8650 519.6000 492.8650 ;
      RECT 506.3000 489.8650 511.4500 492.8650 ;
      RECT 498.1500 489.8650 503.3000 492.8650 ;
      RECT 490.0000 489.8650 495.1500 492.8650 ;
      RECT 481.8500 489.8650 487.0000 492.8650 ;
      RECT 473.7000 489.8650 478.8500 492.8650 ;
      RECT 465.5500 489.8650 470.7000 492.8650 ;
      RECT 457.4000 489.8650 462.5500 492.8650 ;
      RECT 449.2500 489.8650 454.4000 492.8650 ;
      RECT 441.1000 489.8650 446.2500 492.8650 ;
      RECT 432.9500 489.8650 438.1000 492.8650 ;
      RECT 424.8000 489.8650 429.9500 492.8650 ;
      RECT 416.6500 489.8650 421.8000 492.8650 ;
      RECT 396.5000 489.8650 413.6500 492.8650 ;
      RECT 346.5000 489.8650 393.5000 492.8650 ;
      RECT 326.4650 489.8650 343.5000 492.8650 ;
      RECT 317.9500 489.8650 323.4650 492.8650 ;
      RECT 309.4350 489.8650 314.9500 492.8650 ;
      RECT 300.9200 489.8650 306.4350 492.8650 ;
      RECT 292.4050 489.8650 297.9200 492.8650 ;
      RECT 283.8900 489.8650 289.4050 492.8650 ;
      RECT 275.3750 489.8650 280.8900 492.8650 ;
      RECT 266.8600 489.8650 272.3750 492.8650 ;
      RECT 258.3450 489.8650 263.8600 492.8650 ;
      RECT 249.8300 489.8650 255.3450 492.8650 ;
      RECT 241.3150 489.8650 246.8300 492.8650 ;
      RECT 232.8000 489.8650 238.3150 492.8650 ;
      RECT 224.2850 489.8650 229.8000 492.8650 ;
      RECT 215.7700 489.8650 221.2850 492.8650 ;
      RECT 207.2550 489.8650 212.7700 492.8650 ;
      RECT 198.7400 489.8650 204.2550 492.8650 ;
      RECT 190.2250 489.8650 195.7400 492.8650 ;
      RECT 181.7100 489.8650 187.2250 492.8650 ;
      RECT 173.1950 489.8650 178.7100 492.8650 ;
      RECT 164.6800 489.8650 170.1950 492.8650 ;
      RECT 156.1650 489.8650 161.6800 492.8650 ;
      RECT 147.6500 489.8650 153.1650 492.8650 ;
      RECT 139.1350 489.8650 144.6500 492.8650 ;
      RECT 130.6200 489.8650 136.1350 492.8650 ;
      RECT 122.1050 489.8650 127.6200 492.8650 ;
      RECT 113.5900 489.8650 119.1050 492.8650 ;
      RECT 105.0750 489.8650 110.5900 492.8650 ;
      RECT 96.5600 489.8650 102.0750 492.8650 ;
      RECT 88.0450 489.8650 93.5600 492.8650 ;
      RECT 79.5300 489.8650 85.0450 492.8650 ;
      RECT 71.0150 489.8650 76.5300 492.8650 ;
      RECT 62.5000 489.8650 68.0150 492.8650 ;
      RECT 46.5000 489.8650 59.5000 492.8650 ;
      RECT 8.5000 489.8650 43.5000 492.8650 ;
      RECT 0.0000 489.8650 5.5000 492.8650 ;
      RECT 0.0000 488.3000 1120.0000 489.8650 ;
      RECT 1116.6000 487.8650 1120.0000 488.3000 ;
      RECT 0.0000 485.7700 1113.6000 488.3000 ;
      RECT 1118.5000 484.8650 1120.0000 487.8650 ;
      RECT 1114.5000 482.7700 1120.0000 484.8650 ;
      RECT 1076.5000 482.7700 1111.5000 485.7700 ;
      RECT 1060.5000 482.7700 1073.5000 485.7700 ;
      RECT 1052.3500 482.7700 1057.5000 485.7700 ;
      RECT 1044.2000 482.7700 1049.3500 485.7700 ;
      RECT 1036.0500 482.7700 1041.2000 485.7700 ;
      RECT 1027.9000 482.7700 1033.0500 485.7700 ;
      RECT 1019.7500 482.7700 1024.9000 485.7700 ;
      RECT 1011.6000 482.7700 1016.7500 485.7700 ;
      RECT 1003.4500 482.7700 1008.6000 485.7700 ;
      RECT 995.3000 482.7700 1000.4500 485.7700 ;
      RECT 987.1500 482.7700 992.3000 485.7700 ;
      RECT 979.0000 482.7700 984.1500 485.7700 ;
      RECT 970.8500 482.7700 976.0000 485.7700 ;
      RECT 962.7000 482.7700 967.8500 485.7700 ;
      RECT 954.5500 482.7700 959.7000 485.7700 ;
      RECT 946.4000 482.7700 951.5500 485.7700 ;
      RECT 938.2500 482.7700 943.4000 485.7700 ;
      RECT 930.1000 482.7700 935.2500 485.7700 ;
      RECT 921.9500 482.7700 927.1000 485.7700 ;
      RECT 913.8000 482.7700 918.9500 485.7700 ;
      RECT 905.6500 482.7700 910.8000 485.7700 ;
      RECT 897.5000 482.7700 902.6500 485.7700 ;
      RECT 889.3500 482.7700 894.5000 485.7700 ;
      RECT 881.2000 482.7700 886.3500 485.7700 ;
      RECT 873.0500 482.7700 878.2000 485.7700 ;
      RECT 864.9000 482.7700 870.0500 485.7700 ;
      RECT 856.7500 482.7700 861.9000 485.7700 ;
      RECT 848.6000 482.7700 853.7500 485.7700 ;
      RECT 840.4500 482.7700 845.6000 485.7700 ;
      RECT 832.3000 482.7700 837.4500 485.7700 ;
      RECT 824.1500 482.7700 829.3000 485.7700 ;
      RECT 816.0000 482.7700 821.1500 485.7700 ;
      RECT 807.8500 482.7700 813.0000 485.7700 ;
      RECT 799.7000 482.7700 804.8500 485.7700 ;
      RECT 791.5500 482.7700 796.7000 485.7700 ;
      RECT 783.4000 482.7700 788.5500 485.7700 ;
      RECT 775.2500 482.7700 780.4000 485.7700 ;
      RECT 767.1000 482.7700 772.2500 485.7700 ;
      RECT 758.9500 482.7700 764.1000 485.7700 ;
      RECT 750.8000 482.7700 755.9500 485.7700 ;
      RECT 742.6500 482.7700 747.8000 485.7700 ;
      RECT 734.5000 482.7700 739.6500 485.7700 ;
      RECT 726.3500 482.7700 731.5000 485.7700 ;
      RECT 718.2000 482.7700 723.3500 485.7700 ;
      RECT 710.0500 482.7700 715.2000 485.7700 ;
      RECT 701.9000 482.7700 707.0500 485.7700 ;
      RECT 693.7500 482.7700 698.9000 485.7700 ;
      RECT 685.6000 482.7700 690.7500 485.7700 ;
      RECT 677.4500 482.7700 682.6000 485.7700 ;
      RECT 669.3000 482.7700 674.4500 485.7700 ;
      RECT 661.1500 482.7700 666.3000 485.7700 ;
      RECT 653.0000 482.7700 658.1500 485.7700 ;
      RECT 644.8500 482.7700 650.0000 485.7700 ;
      RECT 636.7000 482.7700 641.8500 485.7700 ;
      RECT 628.5500 482.7700 633.7000 485.7700 ;
      RECT 620.4000 482.7700 625.5500 485.7700 ;
      RECT 612.2500 482.7700 617.4000 485.7700 ;
      RECT 604.1000 482.7700 609.2500 485.7700 ;
      RECT 595.9500 482.7700 601.1000 485.7700 ;
      RECT 587.8000 482.7700 592.9500 485.7700 ;
      RECT 579.6500 482.7700 584.8000 485.7700 ;
      RECT 571.5000 482.7700 576.6500 485.7700 ;
      RECT 563.3500 482.7700 568.5000 485.7700 ;
      RECT 555.2000 482.7700 560.3500 485.7700 ;
      RECT 547.0500 482.7700 552.2000 485.7700 ;
      RECT 538.9000 482.7700 544.0500 485.7700 ;
      RECT 530.7500 482.7700 535.9000 485.7700 ;
      RECT 522.6000 482.7700 527.7500 485.7700 ;
      RECT 514.4500 482.7700 519.6000 485.7700 ;
      RECT 506.3000 482.7700 511.4500 485.7700 ;
      RECT 498.1500 482.7700 503.3000 485.7700 ;
      RECT 490.0000 482.7700 495.1500 485.7700 ;
      RECT 481.8500 482.7700 487.0000 485.7700 ;
      RECT 473.7000 482.7700 478.8500 485.7700 ;
      RECT 465.5500 482.7700 470.7000 485.7700 ;
      RECT 457.4000 482.7700 462.5500 485.7700 ;
      RECT 449.2500 482.7700 454.4000 485.7700 ;
      RECT 441.1000 482.7700 446.2500 485.7700 ;
      RECT 432.9500 482.7700 438.1000 485.7700 ;
      RECT 424.8000 482.7700 429.9500 485.7700 ;
      RECT 416.6500 482.7700 421.8000 485.7700 ;
      RECT 396.5000 482.7700 413.6500 485.7700 ;
      RECT 346.5000 482.7700 393.5000 485.7700 ;
      RECT 326.4650 482.7700 343.5000 485.7700 ;
      RECT 317.9500 482.7700 323.4650 485.7700 ;
      RECT 309.4350 482.7700 314.9500 485.7700 ;
      RECT 300.9200 482.7700 306.4350 485.7700 ;
      RECT 292.4050 482.7700 297.9200 485.7700 ;
      RECT 283.8900 482.7700 289.4050 485.7700 ;
      RECT 275.3750 482.7700 280.8900 485.7700 ;
      RECT 266.8600 482.7700 272.3750 485.7700 ;
      RECT 258.3450 482.7700 263.8600 485.7700 ;
      RECT 249.8300 482.7700 255.3450 485.7700 ;
      RECT 241.3150 482.7700 246.8300 485.7700 ;
      RECT 232.8000 482.7700 238.3150 485.7700 ;
      RECT 224.2850 482.7700 229.8000 485.7700 ;
      RECT 215.7700 482.7700 221.2850 485.7700 ;
      RECT 207.2550 482.7700 212.7700 485.7700 ;
      RECT 198.7400 482.7700 204.2550 485.7700 ;
      RECT 190.2250 482.7700 195.7400 485.7700 ;
      RECT 181.7100 482.7700 187.2250 485.7700 ;
      RECT 173.1950 482.7700 178.7100 485.7700 ;
      RECT 164.6800 482.7700 170.1950 485.7700 ;
      RECT 156.1650 482.7700 161.6800 485.7700 ;
      RECT 147.6500 482.7700 153.1650 485.7700 ;
      RECT 139.1350 482.7700 144.6500 485.7700 ;
      RECT 130.6200 482.7700 136.1350 485.7700 ;
      RECT 122.1050 482.7700 127.6200 485.7700 ;
      RECT 113.5900 482.7700 119.1050 485.7700 ;
      RECT 105.0750 482.7700 110.5900 485.7700 ;
      RECT 96.5600 482.7700 102.0750 485.7700 ;
      RECT 88.0450 482.7700 93.5600 485.7700 ;
      RECT 79.5300 482.7700 85.0450 485.7700 ;
      RECT 71.0150 482.7700 76.5300 485.7700 ;
      RECT 62.5000 482.7700 68.0150 485.7700 ;
      RECT 46.5000 482.7700 59.5000 485.7700 ;
      RECT 8.5000 482.7700 43.5000 485.7700 ;
      RECT 0.0000 482.7700 5.5000 485.7700 ;
      RECT 0.0000 481.3000 1120.0000 482.7700 ;
      RECT 1116.6000 480.7700 1120.0000 481.3000 ;
      RECT 0.0000 478.6750 1113.6000 481.3000 ;
      RECT 1118.5000 477.7700 1120.0000 480.7700 ;
      RECT 1114.5000 475.6750 1120.0000 477.7700 ;
      RECT 1076.5000 475.6750 1111.5000 478.6750 ;
      RECT 1060.5000 475.6750 1073.5000 478.6750 ;
      RECT 1052.3500 475.6750 1057.5000 478.6750 ;
      RECT 1044.2000 475.6750 1049.3500 478.6750 ;
      RECT 1036.0500 475.6750 1041.2000 478.6750 ;
      RECT 1027.9000 475.6750 1033.0500 478.6750 ;
      RECT 1019.7500 475.6750 1024.9000 478.6750 ;
      RECT 1011.6000 475.6750 1016.7500 478.6750 ;
      RECT 1003.4500 475.6750 1008.6000 478.6750 ;
      RECT 995.3000 475.6750 1000.4500 478.6750 ;
      RECT 987.1500 475.6750 992.3000 478.6750 ;
      RECT 979.0000 475.6750 984.1500 478.6750 ;
      RECT 970.8500 475.6750 976.0000 478.6750 ;
      RECT 962.7000 475.6750 967.8500 478.6750 ;
      RECT 954.5500 475.6750 959.7000 478.6750 ;
      RECT 946.4000 475.6750 951.5500 478.6750 ;
      RECT 938.2500 475.6750 943.4000 478.6750 ;
      RECT 930.1000 475.6750 935.2500 478.6750 ;
      RECT 921.9500 475.6750 927.1000 478.6750 ;
      RECT 913.8000 475.6750 918.9500 478.6750 ;
      RECT 905.6500 475.6750 910.8000 478.6750 ;
      RECT 897.5000 475.6750 902.6500 478.6750 ;
      RECT 889.3500 475.6750 894.5000 478.6750 ;
      RECT 881.2000 475.6750 886.3500 478.6750 ;
      RECT 873.0500 475.6750 878.2000 478.6750 ;
      RECT 864.9000 475.6750 870.0500 478.6750 ;
      RECT 856.7500 475.6750 861.9000 478.6750 ;
      RECT 848.6000 475.6750 853.7500 478.6750 ;
      RECT 840.4500 475.6750 845.6000 478.6750 ;
      RECT 832.3000 475.6750 837.4500 478.6750 ;
      RECT 824.1500 475.6750 829.3000 478.6750 ;
      RECT 816.0000 475.6750 821.1500 478.6750 ;
      RECT 807.8500 475.6750 813.0000 478.6750 ;
      RECT 799.7000 475.6750 804.8500 478.6750 ;
      RECT 791.5500 475.6750 796.7000 478.6750 ;
      RECT 783.4000 475.6750 788.5500 478.6750 ;
      RECT 775.2500 475.6750 780.4000 478.6750 ;
      RECT 767.1000 475.6750 772.2500 478.6750 ;
      RECT 758.9500 475.6750 764.1000 478.6750 ;
      RECT 750.8000 475.6750 755.9500 478.6750 ;
      RECT 742.6500 475.6750 747.8000 478.6750 ;
      RECT 734.5000 475.6750 739.6500 478.6750 ;
      RECT 726.3500 475.6750 731.5000 478.6750 ;
      RECT 718.2000 475.6750 723.3500 478.6750 ;
      RECT 710.0500 475.6750 715.2000 478.6750 ;
      RECT 701.9000 475.6750 707.0500 478.6750 ;
      RECT 693.7500 475.6750 698.9000 478.6750 ;
      RECT 685.6000 475.6750 690.7500 478.6750 ;
      RECT 677.4500 475.6750 682.6000 478.6750 ;
      RECT 669.3000 475.6750 674.4500 478.6750 ;
      RECT 661.1500 475.6750 666.3000 478.6750 ;
      RECT 653.0000 475.6750 658.1500 478.6750 ;
      RECT 644.8500 475.6750 650.0000 478.6750 ;
      RECT 636.7000 475.6750 641.8500 478.6750 ;
      RECT 628.5500 475.6750 633.7000 478.6750 ;
      RECT 620.4000 475.6750 625.5500 478.6750 ;
      RECT 612.2500 475.6750 617.4000 478.6750 ;
      RECT 604.1000 475.6750 609.2500 478.6750 ;
      RECT 595.9500 475.6750 601.1000 478.6750 ;
      RECT 587.8000 475.6750 592.9500 478.6750 ;
      RECT 579.6500 475.6750 584.8000 478.6750 ;
      RECT 571.5000 475.6750 576.6500 478.6750 ;
      RECT 563.3500 475.6750 568.5000 478.6750 ;
      RECT 555.2000 475.6750 560.3500 478.6750 ;
      RECT 547.0500 475.6750 552.2000 478.6750 ;
      RECT 538.9000 475.6750 544.0500 478.6750 ;
      RECT 530.7500 475.6750 535.9000 478.6750 ;
      RECT 522.6000 475.6750 527.7500 478.6750 ;
      RECT 514.4500 475.6750 519.6000 478.6750 ;
      RECT 506.3000 475.6750 511.4500 478.6750 ;
      RECT 498.1500 475.6750 503.3000 478.6750 ;
      RECT 490.0000 475.6750 495.1500 478.6750 ;
      RECT 481.8500 475.6750 487.0000 478.6750 ;
      RECT 473.7000 475.6750 478.8500 478.6750 ;
      RECT 465.5500 475.6750 470.7000 478.6750 ;
      RECT 457.4000 475.6750 462.5500 478.6750 ;
      RECT 449.2500 475.6750 454.4000 478.6750 ;
      RECT 441.1000 475.6750 446.2500 478.6750 ;
      RECT 432.9500 475.6750 438.1000 478.6750 ;
      RECT 424.8000 475.6750 429.9500 478.6750 ;
      RECT 416.6500 475.6750 421.8000 478.6750 ;
      RECT 396.5000 475.6750 413.6500 478.6750 ;
      RECT 346.5000 475.6750 393.5000 478.6750 ;
      RECT 326.4650 475.6750 343.5000 478.6750 ;
      RECT 317.9500 475.6750 323.4650 478.6750 ;
      RECT 309.4350 475.6750 314.9500 478.6750 ;
      RECT 300.9200 475.6750 306.4350 478.6750 ;
      RECT 292.4050 475.6750 297.9200 478.6750 ;
      RECT 283.8900 475.6750 289.4050 478.6750 ;
      RECT 275.3750 475.6750 280.8900 478.6750 ;
      RECT 266.8600 475.6750 272.3750 478.6750 ;
      RECT 258.3450 475.6750 263.8600 478.6750 ;
      RECT 249.8300 475.6750 255.3450 478.6750 ;
      RECT 241.3150 475.6750 246.8300 478.6750 ;
      RECT 232.8000 475.6750 238.3150 478.6750 ;
      RECT 224.2850 475.6750 229.8000 478.6750 ;
      RECT 215.7700 475.6750 221.2850 478.6750 ;
      RECT 207.2550 475.6750 212.7700 478.6750 ;
      RECT 198.7400 475.6750 204.2550 478.6750 ;
      RECT 190.2250 475.6750 195.7400 478.6750 ;
      RECT 181.7100 475.6750 187.2250 478.6750 ;
      RECT 173.1950 475.6750 178.7100 478.6750 ;
      RECT 164.6800 475.6750 170.1950 478.6750 ;
      RECT 156.1650 475.6750 161.6800 478.6750 ;
      RECT 147.6500 475.6750 153.1650 478.6750 ;
      RECT 139.1350 475.6750 144.6500 478.6750 ;
      RECT 130.6200 475.6750 136.1350 478.6750 ;
      RECT 122.1050 475.6750 127.6200 478.6750 ;
      RECT 113.5900 475.6750 119.1050 478.6750 ;
      RECT 105.0750 475.6750 110.5900 478.6750 ;
      RECT 96.5600 475.6750 102.0750 478.6750 ;
      RECT 88.0450 475.6750 93.5600 478.6750 ;
      RECT 79.5300 475.6750 85.0450 478.6750 ;
      RECT 71.0150 475.6750 76.5300 478.6750 ;
      RECT 62.5000 475.6750 68.0150 478.6750 ;
      RECT 46.5000 475.6750 59.5000 478.6750 ;
      RECT 8.5000 475.6750 43.5000 478.6750 ;
      RECT 0.0000 475.6750 5.5000 478.6750 ;
      RECT 0.0000 474.1000 1120.0000 475.6750 ;
      RECT 1116.6000 473.6750 1120.0000 474.1000 ;
      RECT 0.0000 471.5800 1113.6000 474.1000 ;
      RECT 1118.5000 470.6750 1120.0000 473.6750 ;
      RECT 1114.5000 468.5800 1120.0000 470.6750 ;
      RECT 1076.5000 468.5800 1111.5000 471.5800 ;
      RECT 1060.5000 468.5800 1073.5000 471.5800 ;
      RECT 1052.3500 468.5800 1057.5000 471.5800 ;
      RECT 1044.2000 468.5800 1049.3500 471.5800 ;
      RECT 1036.0500 468.5800 1041.2000 471.5800 ;
      RECT 1027.9000 468.5800 1033.0500 471.5800 ;
      RECT 1019.7500 468.5800 1024.9000 471.5800 ;
      RECT 1011.6000 468.5800 1016.7500 471.5800 ;
      RECT 1003.4500 468.5800 1008.6000 471.5800 ;
      RECT 995.3000 468.5800 1000.4500 471.5800 ;
      RECT 987.1500 468.5800 992.3000 471.5800 ;
      RECT 979.0000 468.5800 984.1500 471.5800 ;
      RECT 970.8500 468.5800 976.0000 471.5800 ;
      RECT 962.7000 468.5800 967.8500 471.5800 ;
      RECT 954.5500 468.5800 959.7000 471.5800 ;
      RECT 946.4000 468.5800 951.5500 471.5800 ;
      RECT 938.2500 468.5800 943.4000 471.5800 ;
      RECT 930.1000 468.5800 935.2500 471.5800 ;
      RECT 921.9500 468.5800 927.1000 471.5800 ;
      RECT 913.8000 468.5800 918.9500 471.5800 ;
      RECT 905.6500 468.5800 910.8000 471.5800 ;
      RECT 897.5000 468.5800 902.6500 471.5800 ;
      RECT 889.3500 468.5800 894.5000 471.5800 ;
      RECT 881.2000 468.5800 886.3500 471.5800 ;
      RECT 873.0500 468.5800 878.2000 471.5800 ;
      RECT 864.9000 468.5800 870.0500 471.5800 ;
      RECT 856.7500 468.5800 861.9000 471.5800 ;
      RECT 848.6000 468.5800 853.7500 471.5800 ;
      RECT 840.4500 468.5800 845.6000 471.5800 ;
      RECT 832.3000 468.5800 837.4500 471.5800 ;
      RECT 824.1500 468.5800 829.3000 471.5800 ;
      RECT 816.0000 468.5800 821.1500 471.5800 ;
      RECT 807.8500 468.5800 813.0000 471.5800 ;
      RECT 799.7000 468.5800 804.8500 471.5800 ;
      RECT 791.5500 468.5800 796.7000 471.5800 ;
      RECT 783.4000 468.5800 788.5500 471.5800 ;
      RECT 775.2500 468.5800 780.4000 471.5800 ;
      RECT 767.1000 468.5800 772.2500 471.5800 ;
      RECT 758.9500 468.5800 764.1000 471.5800 ;
      RECT 750.8000 468.5800 755.9500 471.5800 ;
      RECT 742.6500 468.5800 747.8000 471.5800 ;
      RECT 734.5000 468.5800 739.6500 471.5800 ;
      RECT 726.3500 468.5800 731.5000 471.5800 ;
      RECT 718.2000 468.5800 723.3500 471.5800 ;
      RECT 710.0500 468.5800 715.2000 471.5800 ;
      RECT 701.9000 468.5800 707.0500 471.5800 ;
      RECT 693.7500 468.5800 698.9000 471.5800 ;
      RECT 685.6000 468.5800 690.7500 471.5800 ;
      RECT 677.4500 468.5800 682.6000 471.5800 ;
      RECT 669.3000 468.5800 674.4500 471.5800 ;
      RECT 661.1500 468.5800 666.3000 471.5800 ;
      RECT 653.0000 468.5800 658.1500 471.5800 ;
      RECT 644.8500 468.5800 650.0000 471.5800 ;
      RECT 636.7000 468.5800 641.8500 471.5800 ;
      RECT 628.5500 468.5800 633.7000 471.5800 ;
      RECT 620.4000 468.5800 625.5500 471.5800 ;
      RECT 612.2500 468.5800 617.4000 471.5800 ;
      RECT 604.1000 468.5800 609.2500 471.5800 ;
      RECT 595.9500 468.5800 601.1000 471.5800 ;
      RECT 587.8000 468.5800 592.9500 471.5800 ;
      RECT 579.6500 468.5800 584.8000 471.5800 ;
      RECT 571.5000 468.5800 576.6500 471.5800 ;
      RECT 563.3500 468.5800 568.5000 471.5800 ;
      RECT 555.2000 468.5800 560.3500 471.5800 ;
      RECT 547.0500 468.5800 552.2000 471.5800 ;
      RECT 538.9000 468.5800 544.0500 471.5800 ;
      RECT 530.7500 468.5800 535.9000 471.5800 ;
      RECT 522.6000 468.5800 527.7500 471.5800 ;
      RECT 514.4500 468.5800 519.6000 471.5800 ;
      RECT 506.3000 468.5800 511.4500 471.5800 ;
      RECT 498.1500 468.5800 503.3000 471.5800 ;
      RECT 490.0000 468.5800 495.1500 471.5800 ;
      RECT 481.8500 468.5800 487.0000 471.5800 ;
      RECT 473.7000 468.5800 478.8500 471.5800 ;
      RECT 465.5500 468.5800 470.7000 471.5800 ;
      RECT 457.4000 468.5800 462.5500 471.5800 ;
      RECT 449.2500 468.5800 454.4000 471.5800 ;
      RECT 441.1000 468.5800 446.2500 471.5800 ;
      RECT 432.9500 468.5800 438.1000 471.5800 ;
      RECT 424.8000 468.5800 429.9500 471.5800 ;
      RECT 416.6500 468.5800 421.8000 471.5800 ;
      RECT 396.5000 468.5800 413.6500 471.5800 ;
      RECT 346.5000 468.5800 393.5000 471.5800 ;
      RECT 326.4650 468.5800 343.5000 471.5800 ;
      RECT 317.9500 468.5800 323.4650 471.5800 ;
      RECT 309.4350 468.5800 314.9500 471.5800 ;
      RECT 300.9200 468.5800 306.4350 471.5800 ;
      RECT 292.4050 468.5800 297.9200 471.5800 ;
      RECT 283.8900 468.5800 289.4050 471.5800 ;
      RECT 275.3750 468.5800 280.8900 471.5800 ;
      RECT 266.8600 468.5800 272.3750 471.5800 ;
      RECT 258.3450 468.5800 263.8600 471.5800 ;
      RECT 249.8300 468.5800 255.3450 471.5800 ;
      RECT 241.3150 468.5800 246.8300 471.5800 ;
      RECT 232.8000 468.5800 238.3150 471.5800 ;
      RECT 224.2850 468.5800 229.8000 471.5800 ;
      RECT 215.7700 468.5800 221.2850 471.5800 ;
      RECT 207.2550 468.5800 212.7700 471.5800 ;
      RECT 198.7400 468.5800 204.2550 471.5800 ;
      RECT 190.2250 468.5800 195.7400 471.5800 ;
      RECT 181.7100 468.5800 187.2250 471.5800 ;
      RECT 173.1950 468.5800 178.7100 471.5800 ;
      RECT 164.6800 468.5800 170.1950 471.5800 ;
      RECT 156.1650 468.5800 161.6800 471.5800 ;
      RECT 147.6500 468.5800 153.1650 471.5800 ;
      RECT 139.1350 468.5800 144.6500 471.5800 ;
      RECT 130.6200 468.5800 136.1350 471.5800 ;
      RECT 122.1050 468.5800 127.6200 471.5800 ;
      RECT 113.5900 468.5800 119.1050 471.5800 ;
      RECT 105.0750 468.5800 110.5900 471.5800 ;
      RECT 96.5600 468.5800 102.0750 471.5800 ;
      RECT 88.0450 468.5800 93.5600 471.5800 ;
      RECT 79.5300 468.5800 85.0450 471.5800 ;
      RECT 71.0150 468.5800 76.5300 471.5800 ;
      RECT 62.5000 468.5800 68.0150 471.5800 ;
      RECT 46.5000 468.5800 59.5000 471.5800 ;
      RECT 8.5000 468.5800 43.5000 471.5800 ;
      RECT 0.0000 468.5800 5.5000 471.5800 ;
      RECT 0.0000 467.1000 1120.0000 468.5800 ;
      RECT 1116.6000 466.5800 1120.0000 467.1000 ;
      RECT 0.0000 464.4850 1113.6000 467.1000 ;
      RECT 1118.5000 463.5800 1120.0000 466.5800 ;
      RECT 1114.5000 461.4850 1120.0000 463.5800 ;
      RECT 1076.5000 461.4850 1111.5000 464.4850 ;
      RECT 1060.5000 461.4850 1073.5000 464.4850 ;
      RECT 1052.3500 461.4850 1057.5000 464.4850 ;
      RECT 1044.2000 461.4850 1049.3500 464.4850 ;
      RECT 1036.0500 461.4850 1041.2000 464.4850 ;
      RECT 1027.9000 461.4850 1033.0500 464.4850 ;
      RECT 1019.7500 461.4850 1024.9000 464.4850 ;
      RECT 1011.6000 461.4850 1016.7500 464.4850 ;
      RECT 1003.4500 461.4850 1008.6000 464.4850 ;
      RECT 995.3000 461.4850 1000.4500 464.4850 ;
      RECT 987.1500 461.4850 992.3000 464.4850 ;
      RECT 979.0000 461.4850 984.1500 464.4850 ;
      RECT 970.8500 461.4850 976.0000 464.4850 ;
      RECT 962.7000 461.4850 967.8500 464.4850 ;
      RECT 954.5500 461.4850 959.7000 464.4850 ;
      RECT 946.4000 461.4850 951.5500 464.4850 ;
      RECT 938.2500 461.4850 943.4000 464.4850 ;
      RECT 930.1000 461.4850 935.2500 464.4850 ;
      RECT 921.9500 461.4850 927.1000 464.4850 ;
      RECT 913.8000 461.4850 918.9500 464.4850 ;
      RECT 905.6500 461.4850 910.8000 464.4850 ;
      RECT 897.5000 461.4850 902.6500 464.4850 ;
      RECT 889.3500 461.4850 894.5000 464.4850 ;
      RECT 881.2000 461.4850 886.3500 464.4850 ;
      RECT 873.0500 461.4850 878.2000 464.4850 ;
      RECT 864.9000 461.4850 870.0500 464.4850 ;
      RECT 856.7500 461.4850 861.9000 464.4850 ;
      RECT 848.6000 461.4850 853.7500 464.4850 ;
      RECT 840.4500 461.4850 845.6000 464.4850 ;
      RECT 832.3000 461.4850 837.4500 464.4850 ;
      RECT 824.1500 461.4850 829.3000 464.4850 ;
      RECT 816.0000 461.4850 821.1500 464.4850 ;
      RECT 807.8500 461.4850 813.0000 464.4850 ;
      RECT 799.7000 461.4850 804.8500 464.4850 ;
      RECT 791.5500 461.4850 796.7000 464.4850 ;
      RECT 783.4000 461.4850 788.5500 464.4850 ;
      RECT 775.2500 461.4850 780.4000 464.4850 ;
      RECT 767.1000 461.4850 772.2500 464.4850 ;
      RECT 758.9500 461.4850 764.1000 464.4850 ;
      RECT 750.8000 461.4850 755.9500 464.4850 ;
      RECT 742.6500 461.4850 747.8000 464.4850 ;
      RECT 734.5000 461.4850 739.6500 464.4850 ;
      RECT 726.3500 461.4850 731.5000 464.4850 ;
      RECT 718.2000 461.4850 723.3500 464.4850 ;
      RECT 710.0500 461.4850 715.2000 464.4850 ;
      RECT 701.9000 461.4850 707.0500 464.4850 ;
      RECT 693.7500 461.4850 698.9000 464.4850 ;
      RECT 685.6000 461.4850 690.7500 464.4850 ;
      RECT 677.4500 461.4850 682.6000 464.4850 ;
      RECT 669.3000 461.4850 674.4500 464.4850 ;
      RECT 661.1500 461.4850 666.3000 464.4850 ;
      RECT 653.0000 461.4850 658.1500 464.4850 ;
      RECT 644.8500 461.4850 650.0000 464.4850 ;
      RECT 636.7000 461.4850 641.8500 464.4850 ;
      RECT 628.5500 461.4850 633.7000 464.4850 ;
      RECT 620.4000 461.4850 625.5500 464.4850 ;
      RECT 612.2500 461.4850 617.4000 464.4850 ;
      RECT 604.1000 461.4850 609.2500 464.4850 ;
      RECT 595.9500 461.4850 601.1000 464.4850 ;
      RECT 587.8000 461.4850 592.9500 464.4850 ;
      RECT 579.6500 461.4850 584.8000 464.4850 ;
      RECT 571.5000 461.4850 576.6500 464.4850 ;
      RECT 563.3500 461.4850 568.5000 464.4850 ;
      RECT 555.2000 461.4850 560.3500 464.4850 ;
      RECT 547.0500 461.4850 552.2000 464.4850 ;
      RECT 538.9000 461.4850 544.0500 464.4850 ;
      RECT 530.7500 461.4850 535.9000 464.4850 ;
      RECT 522.6000 461.4850 527.7500 464.4850 ;
      RECT 514.4500 461.4850 519.6000 464.4850 ;
      RECT 506.3000 461.4850 511.4500 464.4850 ;
      RECT 498.1500 461.4850 503.3000 464.4850 ;
      RECT 490.0000 461.4850 495.1500 464.4850 ;
      RECT 481.8500 461.4850 487.0000 464.4850 ;
      RECT 473.7000 461.4850 478.8500 464.4850 ;
      RECT 465.5500 461.4850 470.7000 464.4850 ;
      RECT 457.4000 461.4850 462.5500 464.4850 ;
      RECT 449.2500 461.4850 454.4000 464.4850 ;
      RECT 441.1000 461.4850 446.2500 464.4850 ;
      RECT 432.9500 461.4850 438.1000 464.4850 ;
      RECT 424.8000 461.4850 429.9500 464.4850 ;
      RECT 416.6500 461.4850 421.8000 464.4850 ;
      RECT 396.5000 461.4850 413.6500 464.4850 ;
      RECT 346.5000 461.4850 393.5000 464.4850 ;
      RECT 326.4650 461.4850 343.5000 464.4850 ;
      RECT 317.9500 461.4850 323.4650 464.4850 ;
      RECT 309.4350 461.4850 314.9500 464.4850 ;
      RECT 300.9200 461.4850 306.4350 464.4850 ;
      RECT 292.4050 461.4850 297.9200 464.4850 ;
      RECT 283.8900 461.4850 289.4050 464.4850 ;
      RECT 275.3750 461.4850 280.8900 464.4850 ;
      RECT 266.8600 461.4850 272.3750 464.4850 ;
      RECT 258.3450 461.4850 263.8600 464.4850 ;
      RECT 249.8300 461.4850 255.3450 464.4850 ;
      RECT 241.3150 461.4850 246.8300 464.4850 ;
      RECT 232.8000 461.4850 238.3150 464.4850 ;
      RECT 224.2850 461.4850 229.8000 464.4850 ;
      RECT 215.7700 461.4850 221.2850 464.4850 ;
      RECT 207.2550 461.4850 212.7700 464.4850 ;
      RECT 198.7400 461.4850 204.2550 464.4850 ;
      RECT 190.2250 461.4850 195.7400 464.4850 ;
      RECT 181.7100 461.4850 187.2250 464.4850 ;
      RECT 173.1950 461.4850 178.7100 464.4850 ;
      RECT 164.6800 461.4850 170.1950 464.4850 ;
      RECT 156.1650 461.4850 161.6800 464.4850 ;
      RECT 147.6500 461.4850 153.1650 464.4850 ;
      RECT 139.1350 461.4850 144.6500 464.4850 ;
      RECT 130.6200 461.4850 136.1350 464.4850 ;
      RECT 122.1050 461.4850 127.6200 464.4850 ;
      RECT 113.5900 461.4850 119.1050 464.4850 ;
      RECT 105.0750 461.4850 110.5900 464.4850 ;
      RECT 96.5600 461.4850 102.0750 464.4850 ;
      RECT 88.0450 461.4850 93.5600 464.4850 ;
      RECT 79.5300 461.4850 85.0450 464.4850 ;
      RECT 71.0150 461.4850 76.5300 464.4850 ;
      RECT 62.5000 461.4850 68.0150 464.4850 ;
      RECT 46.5000 461.4850 59.5000 464.4850 ;
      RECT 8.5000 461.4850 43.5000 464.4850 ;
      RECT 0.0000 461.4850 5.5000 464.4850 ;
      RECT 0.0000 459.9000 1120.0000 461.4850 ;
      RECT 1116.6000 459.4850 1120.0000 459.9000 ;
      RECT 0.0000 457.3900 1113.6000 459.9000 ;
      RECT 1118.5000 456.4850 1120.0000 459.4850 ;
      RECT 1114.5000 454.3900 1120.0000 456.4850 ;
      RECT 1076.5000 454.3900 1111.5000 457.3900 ;
      RECT 1060.5000 454.3900 1073.5000 457.3900 ;
      RECT 1052.3500 454.3900 1057.5000 457.3900 ;
      RECT 1044.2000 454.3900 1049.3500 457.3900 ;
      RECT 1036.0500 454.3900 1041.2000 457.3900 ;
      RECT 1027.9000 454.3900 1033.0500 457.3900 ;
      RECT 1019.7500 454.3900 1024.9000 457.3900 ;
      RECT 1011.6000 454.3900 1016.7500 457.3900 ;
      RECT 1003.4500 454.3900 1008.6000 457.3900 ;
      RECT 995.3000 454.3900 1000.4500 457.3900 ;
      RECT 987.1500 454.3900 992.3000 457.3900 ;
      RECT 979.0000 454.3900 984.1500 457.3900 ;
      RECT 970.8500 454.3900 976.0000 457.3900 ;
      RECT 962.7000 454.3900 967.8500 457.3900 ;
      RECT 954.5500 454.3900 959.7000 457.3900 ;
      RECT 946.4000 454.3900 951.5500 457.3900 ;
      RECT 938.2500 454.3900 943.4000 457.3900 ;
      RECT 930.1000 454.3900 935.2500 457.3900 ;
      RECT 921.9500 454.3900 927.1000 457.3900 ;
      RECT 913.8000 454.3900 918.9500 457.3900 ;
      RECT 905.6500 454.3900 910.8000 457.3900 ;
      RECT 897.5000 454.3900 902.6500 457.3900 ;
      RECT 889.3500 454.3900 894.5000 457.3900 ;
      RECT 881.2000 454.3900 886.3500 457.3900 ;
      RECT 873.0500 454.3900 878.2000 457.3900 ;
      RECT 864.9000 454.3900 870.0500 457.3900 ;
      RECT 856.7500 454.3900 861.9000 457.3900 ;
      RECT 848.6000 454.3900 853.7500 457.3900 ;
      RECT 840.4500 454.3900 845.6000 457.3900 ;
      RECT 832.3000 454.3900 837.4500 457.3900 ;
      RECT 824.1500 454.3900 829.3000 457.3900 ;
      RECT 816.0000 454.3900 821.1500 457.3900 ;
      RECT 807.8500 454.3900 813.0000 457.3900 ;
      RECT 799.7000 454.3900 804.8500 457.3900 ;
      RECT 791.5500 454.3900 796.7000 457.3900 ;
      RECT 783.4000 454.3900 788.5500 457.3900 ;
      RECT 775.2500 454.3900 780.4000 457.3900 ;
      RECT 767.1000 454.3900 772.2500 457.3900 ;
      RECT 758.9500 454.3900 764.1000 457.3900 ;
      RECT 750.8000 454.3900 755.9500 457.3900 ;
      RECT 742.6500 454.3900 747.8000 457.3900 ;
      RECT 734.5000 454.3900 739.6500 457.3900 ;
      RECT 726.3500 454.3900 731.5000 457.3900 ;
      RECT 718.2000 454.3900 723.3500 457.3900 ;
      RECT 710.0500 454.3900 715.2000 457.3900 ;
      RECT 701.9000 454.3900 707.0500 457.3900 ;
      RECT 693.7500 454.3900 698.9000 457.3900 ;
      RECT 685.6000 454.3900 690.7500 457.3900 ;
      RECT 677.4500 454.3900 682.6000 457.3900 ;
      RECT 669.3000 454.3900 674.4500 457.3900 ;
      RECT 661.1500 454.3900 666.3000 457.3900 ;
      RECT 653.0000 454.3900 658.1500 457.3900 ;
      RECT 644.8500 454.3900 650.0000 457.3900 ;
      RECT 636.7000 454.3900 641.8500 457.3900 ;
      RECT 628.5500 454.3900 633.7000 457.3900 ;
      RECT 620.4000 454.3900 625.5500 457.3900 ;
      RECT 612.2500 454.3900 617.4000 457.3900 ;
      RECT 604.1000 454.3900 609.2500 457.3900 ;
      RECT 595.9500 454.3900 601.1000 457.3900 ;
      RECT 587.8000 454.3900 592.9500 457.3900 ;
      RECT 579.6500 454.3900 584.8000 457.3900 ;
      RECT 571.5000 454.3900 576.6500 457.3900 ;
      RECT 563.3500 454.3900 568.5000 457.3900 ;
      RECT 555.2000 454.3900 560.3500 457.3900 ;
      RECT 547.0500 454.3900 552.2000 457.3900 ;
      RECT 538.9000 454.3900 544.0500 457.3900 ;
      RECT 530.7500 454.3900 535.9000 457.3900 ;
      RECT 522.6000 454.3900 527.7500 457.3900 ;
      RECT 514.4500 454.3900 519.6000 457.3900 ;
      RECT 506.3000 454.3900 511.4500 457.3900 ;
      RECT 498.1500 454.3900 503.3000 457.3900 ;
      RECT 490.0000 454.3900 495.1500 457.3900 ;
      RECT 481.8500 454.3900 487.0000 457.3900 ;
      RECT 473.7000 454.3900 478.8500 457.3900 ;
      RECT 465.5500 454.3900 470.7000 457.3900 ;
      RECT 457.4000 454.3900 462.5500 457.3900 ;
      RECT 449.2500 454.3900 454.4000 457.3900 ;
      RECT 441.1000 454.3900 446.2500 457.3900 ;
      RECT 432.9500 454.3900 438.1000 457.3900 ;
      RECT 424.8000 454.3900 429.9500 457.3900 ;
      RECT 416.6500 454.3900 421.8000 457.3900 ;
      RECT 396.5000 454.3900 413.6500 457.3900 ;
      RECT 346.5000 454.3900 393.5000 457.3900 ;
      RECT 326.4650 454.3900 343.5000 457.3900 ;
      RECT 317.9500 454.3900 323.4650 457.3900 ;
      RECT 309.4350 454.3900 314.9500 457.3900 ;
      RECT 300.9200 454.3900 306.4350 457.3900 ;
      RECT 292.4050 454.3900 297.9200 457.3900 ;
      RECT 283.8900 454.3900 289.4050 457.3900 ;
      RECT 275.3750 454.3900 280.8900 457.3900 ;
      RECT 266.8600 454.3900 272.3750 457.3900 ;
      RECT 258.3450 454.3900 263.8600 457.3900 ;
      RECT 249.8300 454.3900 255.3450 457.3900 ;
      RECT 241.3150 454.3900 246.8300 457.3900 ;
      RECT 232.8000 454.3900 238.3150 457.3900 ;
      RECT 224.2850 454.3900 229.8000 457.3900 ;
      RECT 215.7700 454.3900 221.2850 457.3900 ;
      RECT 207.2550 454.3900 212.7700 457.3900 ;
      RECT 198.7400 454.3900 204.2550 457.3900 ;
      RECT 190.2250 454.3900 195.7400 457.3900 ;
      RECT 181.7100 454.3900 187.2250 457.3900 ;
      RECT 173.1950 454.3900 178.7100 457.3900 ;
      RECT 164.6800 454.3900 170.1950 457.3900 ;
      RECT 156.1650 454.3900 161.6800 457.3900 ;
      RECT 147.6500 454.3900 153.1650 457.3900 ;
      RECT 139.1350 454.3900 144.6500 457.3900 ;
      RECT 130.6200 454.3900 136.1350 457.3900 ;
      RECT 122.1050 454.3900 127.6200 457.3900 ;
      RECT 113.5900 454.3900 119.1050 457.3900 ;
      RECT 105.0750 454.3900 110.5900 457.3900 ;
      RECT 96.5600 454.3900 102.0750 457.3900 ;
      RECT 88.0450 454.3900 93.5600 457.3900 ;
      RECT 79.5300 454.3900 85.0450 457.3900 ;
      RECT 71.0150 454.3900 76.5300 457.3900 ;
      RECT 62.5000 454.3900 68.0150 457.3900 ;
      RECT 46.5000 454.3900 59.5000 457.3900 ;
      RECT 8.5000 454.3900 43.5000 457.3900 ;
      RECT 0.0000 454.3900 5.5000 457.3900 ;
      RECT 0.0000 452.9000 1120.0000 454.3900 ;
      RECT 1116.6000 452.3900 1120.0000 452.9000 ;
      RECT 0.0000 450.2950 1113.6000 452.9000 ;
      RECT 1118.5000 449.3900 1120.0000 452.3900 ;
      RECT 1114.5000 447.2950 1120.0000 449.3900 ;
      RECT 1076.5000 447.2950 1111.5000 450.2950 ;
      RECT 1060.5000 447.2950 1073.5000 450.2950 ;
      RECT 1052.3500 447.2950 1057.5000 450.2950 ;
      RECT 1044.2000 447.2950 1049.3500 450.2950 ;
      RECT 1036.0500 447.2950 1041.2000 450.2950 ;
      RECT 1027.9000 447.2950 1033.0500 450.2950 ;
      RECT 1019.7500 447.2950 1024.9000 450.2950 ;
      RECT 1011.6000 447.2950 1016.7500 450.2950 ;
      RECT 1003.4500 447.2950 1008.6000 450.2950 ;
      RECT 995.3000 447.2950 1000.4500 450.2950 ;
      RECT 987.1500 447.2950 992.3000 450.2950 ;
      RECT 979.0000 447.2950 984.1500 450.2950 ;
      RECT 970.8500 447.2950 976.0000 450.2950 ;
      RECT 962.7000 447.2950 967.8500 450.2950 ;
      RECT 954.5500 447.2950 959.7000 450.2950 ;
      RECT 946.4000 447.2950 951.5500 450.2950 ;
      RECT 938.2500 447.2950 943.4000 450.2950 ;
      RECT 930.1000 447.2950 935.2500 450.2950 ;
      RECT 921.9500 447.2950 927.1000 450.2950 ;
      RECT 913.8000 447.2950 918.9500 450.2950 ;
      RECT 905.6500 447.2950 910.8000 450.2950 ;
      RECT 897.5000 447.2950 902.6500 450.2950 ;
      RECT 889.3500 447.2950 894.5000 450.2950 ;
      RECT 881.2000 447.2950 886.3500 450.2950 ;
      RECT 873.0500 447.2950 878.2000 450.2950 ;
      RECT 864.9000 447.2950 870.0500 450.2950 ;
      RECT 856.7500 447.2950 861.9000 450.2950 ;
      RECT 848.6000 447.2950 853.7500 450.2950 ;
      RECT 840.4500 447.2950 845.6000 450.2950 ;
      RECT 832.3000 447.2950 837.4500 450.2950 ;
      RECT 824.1500 447.2950 829.3000 450.2950 ;
      RECT 816.0000 447.2950 821.1500 450.2950 ;
      RECT 807.8500 447.2950 813.0000 450.2950 ;
      RECT 799.7000 447.2950 804.8500 450.2950 ;
      RECT 791.5500 447.2950 796.7000 450.2950 ;
      RECT 783.4000 447.2950 788.5500 450.2950 ;
      RECT 775.2500 447.2950 780.4000 450.2950 ;
      RECT 767.1000 447.2950 772.2500 450.2950 ;
      RECT 758.9500 447.2950 764.1000 450.2950 ;
      RECT 750.8000 447.2950 755.9500 450.2950 ;
      RECT 742.6500 447.2950 747.8000 450.2950 ;
      RECT 734.5000 447.2950 739.6500 450.2950 ;
      RECT 726.3500 447.2950 731.5000 450.2950 ;
      RECT 718.2000 447.2950 723.3500 450.2950 ;
      RECT 710.0500 447.2950 715.2000 450.2950 ;
      RECT 701.9000 447.2950 707.0500 450.2950 ;
      RECT 693.7500 447.2950 698.9000 450.2950 ;
      RECT 685.6000 447.2950 690.7500 450.2950 ;
      RECT 677.4500 447.2950 682.6000 450.2950 ;
      RECT 669.3000 447.2950 674.4500 450.2950 ;
      RECT 661.1500 447.2950 666.3000 450.2950 ;
      RECT 653.0000 447.2950 658.1500 450.2950 ;
      RECT 644.8500 447.2950 650.0000 450.2950 ;
      RECT 636.7000 447.2950 641.8500 450.2950 ;
      RECT 628.5500 447.2950 633.7000 450.2950 ;
      RECT 620.4000 447.2950 625.5500 450.2950 ;
      RECT 612.2500 447.2950 617.4000 450.2950 ;
      RECT 604.1000 447.2950 609.2500 450.2950 ;
      RECT 595.9500 447.2950 601.1000 450.2950 ;
      RECT 587.8000 447.2950 592.9500 450.2950 ;
      RECT 579.6500 447.2950 584.8000 450.2950 ;
      RECT 571.5000 447.2950 576.6500 450.2950 ;
      RECT 563.3500 447.2950 568.5000 450.2950 ;
      RECT 555.2000 447.2950 560.3500 450.2950 ;
      RECT 547.0500 447.2950 552.2000 450.2950 ;
      RECT 538.9000 447.2950 544.0500 450.2950 ;
      RECT 530.7500 447.2950 535.9000 450.2950 ;
      RECT 522.6000 447.2950 527.7500 450.2950 ;
      RECT 514.4500 447.2950 519.6000 450.2950 ;
      RECT 506.3000 447.2950 511.4500 450.2950 ;
      RECT 498.1500 447.2950 503.3000 450.2950 ;
      RECT 490.0000 447.2950 495.1500 450.2950 ;
      RECT 481.8500 447.2950 487.0000 450.2950 ;
      RECT 473.7000 447.2950 478.8500 450.2950 ;
      RECT 465.5500 447.2950 470.7000 450.2950 ;
      RECT 457.4000 447.2950 462.5500 450.2950 ;
      RECT 449.2500 447.2950 454.4000 450.2950 ;
      RECT 441.1000 447.2950 446.2500 450.2950 ;
      RECT 432.9500 447.2950 438.1000 450.2950 ;
      RECT 424.8000 447.2950 429.9500 450.2950 ;
      RECT 416.6500 447.2950 421.8000 450.2950 ;
      RECT 396.5000 447.2950 413.6500 450.2950 ;
      RECT 346.5000 447.2950 393.5000 450.2950 ;
      RECT 326.4650 447.2950 343.5000 450.2950 ;
      RECT 317.9500 447.2950 323.4650 450.2950 ;
      RECT 309.4350 447.2950 314.9500 450.2950 ;
      RECT 300.9200 447.2950 306.4350 450.2950 ;
      RECT 292.4050 447.2950 297.9200 450.2950 ;
      RECT 283.8900 447.2950 289.4050 450.2950 ;
      RECT 275.3750 447.2950 280.8900 450.2950 ;
      RECT 266.8600 447.2950 272.3750 450.2950 ;
      RECT 258.3450 447.2950 263.8600 450.2950 ;
      RECT 249.8300 447.2950 255.3450 450.2950 ;
      RECT 241.3150 447.2950 246.8300 450.2950 ;
      RECT 232.8000 447.2950 238.3150 450.2950 ;
      RECT 224.2850 447.2950 229.8000 450.2950 ;
      RECT 215.7700 447.2950 221.2850 450.2950 ;
      RECT 207.2550 447.2950 212.7700 450.2950 ;
      RECT 198.7400 447.2950 204.2550 450.2950 ;
      RECT 190.2250 447.2950 195.7400 450.2950 ;
      RECT 181.7100 447.2950 187.2250 450.2950 ;
      RECT 173.1950 447.2950 178.7100 450.2950 ;
      RECT 164.6800 447.2950 170.1950 450.2950 ;
      RECT 156.1650 447.2950 161.6800 450.2950 ;
      RECT 147.6500 447.2950 153.1650 450.2950 ;
      RECT 139.1350 447.2950 144.6500 450.2950 ;
      RECT 130.6200 447.2950 136.1350 450.2950 ;
      RECT 122.1050 447.2950 127.6200 450.2950 ;
      RECT 113.5900 447.2950 119.1050 450.2950 ;
      RECT 105.0750 447.2950 110.5900 450.2950 ;
      RECT 96.5600 447.2950 102.0750 450.2950 ;
      RECT 88.0450 447.2950 93.5600 450.2950 ;
      RECT 79.5300 447.2950 85.0450 450.2950 ;
      RECT 71.0150 447.2950 76.5300 450.2950 ;
      RECT 62.5000 447.2950 68.0150 450.2950 ;
      RECT 46.5000 447.2950 59.5000 450.2950 ;
      RECT 8.5000 447.2950 43.5000 450.2950 ;
      RECT 0.0000 447.2950 5.5000 450.2950 ;
      RECT 0.0000 445.7000 1120.0000 447.2950 ;
      RECT 1116.6000 445.2950 1120.0000 445.7000 ;
      RECT 0.0000 443.2000 1113.6000 445.7000 ;
      RECT 1118.5000 442.2950 1120.0000 445.2950 ;
      RECT 1114.5000 440.2000 1120.0000 442.2950 ;
      RECT 1076.5000 440.2000 1111.5000 443.2000 ;
      RECT 1060.5000 440.2000 1073.5000 443.2000 ;
      RECT 1052.3500 440.2000 1057.5000 443.2000 ;
      RECT 1044.2000 440.2000 1049.3500 443.2000 ;
      RECT 1036.0500 440.2000 1041.2000 443.2000 ;
      RECT 1027.9000 440.2000 1033.0500 443.2000 ;
      RECT 1019.7500 440.2000 1024.9000 443.2000 ;
      RECT 1011.6000 440.2000 1016.7500 443.2000 ;
      RECT 1003.4500 440.2000 1008.6000 443.2000 ;
      RECT 995.3000 440.2000 1000.4500 443.2000 ;
      RECT 987.1500 440.2000 992.3000 443.2000 ;
      RECT 979.0000 440.2000 984.1500 443.2000 ;
      RECT 970.8500 440.2000 976.0000 443.2000 ;
      RECT 962.7000 440.2000 967.8500 443.2000 ;
      RECT 954.5500 440.2000 959.7000 443.2000 ;
      RECT 946.4000 440.2000 951.5500 443.2000 ;
      RECT 938.2500 440.2000 943.4000 443.2000 ;
      RECT 930.1000 440.2000 935.2500 443.2000 ;
      RECT 921.9500 440.2000 927.1000 443.2000 ;
      RECT 913.8000 440.2000 918.9500 443.2000 ;
      RECT 905.6500 440.2000 910.8000 443.2000 ;
      RECT 897.5000 440.2000 902.6500 443.2000 ;
      RECT 889.3500 440.2000 894.5000 443.2000 ;
      RECT 881.2000 440.2000 886.3500 443.2000 ;
      RECT 873.0500 440.2000 878.2000 443.2000 ;
      RECT 864.9000 440.2000 870.0500 443.2000 ;
      RECT 856.7500 440.2000 861.9000 443.2000 ;
      RECT 848.6000 440.2000 853.7500 443.2000 ;
      RECT 840.4500 440.2000 845.6000 443.2000 ;
      RECT 832.3000 440.2000 837.4500 443.2000 ;
      RECT 824.1500 440.2000 829.3000 443.2000 ;
      RECT 816.0000 440.2000 821.1500 443.2000 ;
      RECT 807.8500 440.2000 813.0000 443.2000 ;
      RECT 799.7000 440.2000 804.8500 443.2000 ;
      RECT 791.5500 440.2000 796.7000 443.2000 ;
      RECT 783.4000 440.2000 788.5500 443.2000 ;
      RECT 775.2500 440.2000 780.4000 443.2000 ;
      RECT 767.1000 440.2000 772.2500 443.2000 ;
      RECT 758.9500 440.2000 764.1000 443.2000 ;
      RECT 750.8000 440.2000 755.9500 443.2000 ;
      RECT 742.6500 440.2000 747.8000 443.2000 ;
      RECT 734.5000 440.2000 739.6500 443.2000 ;
      RECT 726.3500 440.2000 731.5000 443.2000 ;
      RECT 718.2000 440.2000 723.3500 443.2000 ;
      RECT 710.0500 440.2000 715.2000 443.2000 ;
      RECT 701.9000 440.2000 707.0500 443.2000 ;
      RECT 693.7500 440.2000 698.9000 443.2000 ;
      RECT 685.6000 440.2000 690.7500 443.2000 ;
      RECT 677.4500 440.2000 682.6000 443.2000 ;
      RECT 669.3000 440.2000 674.4500 443.2000 ;
      RECT 661.1500 440.2000 666.3000 443.2000 ;
      RECT 653.0000 440.2000 658.1500 443.2000 ;
      RECT 644.8500 440.2000 650.0000 443.2000 ;
      RECT 636.7000 440.2000 641.8500 443.2000 ;
      RECT 628.5500 440.2000 633.7000 443.2000 ;
      RECT 620.4000 440.2000 625.5500 443.2000 ;
      RECT 612.2500 440.2000 617.4000 443.2000 ;
      RECT 604.1000 440.2000 609.2500 443.2000 ;
      RECT 595.9500 440.2000 601.1000 443.2000 ;
      RECT 587.8000 440.2000 592.9500 443.2000 ;
      RECT 579.6500 440.2000 584.8000 443.2000 ;
      RECT 571.5000 440.2000 576.6500 443.2000 ;
      RECT 563.3500 440.2000 568.5000 443.2000 ;
      RECT 555.2000 440.2000 560.3500 443.2000 ;
      RECT 547.0500 440.2000 552.2000 443.2000 ;
      RECT 538.9000 440.2000 544.0500 443.2000 ;
      RECT 530.7500 440.2000 535.9000 443.2000 ;
      RECT 522.6000 440.2000 527.7500 443.2000 ;
      RECT 514.4500 440.2000 519.6000 443.2000 ;
      RECT 506.3000 440.2000 511.4500 443.2000 ;
      RECT 498.1500 440.2000 503.3000 443.2000 ;
      RECT 490.0000 440.2000 495.1500 443.2000 ;
      RECT 481.8500 440.2000 487.0000 443.2000 ;
      RECT 473.7000 440.2000 478.8500 443.2000 ;
      RECT 465.5500 440.2000 470.7000 443.2000 ;
      RECT 457.4000 440.2000 462.5500 443.2000 ;
      RECT 449.2500 440.2000 454.4000 443.2000 ;
      RECT 441.1000 440.2000 446.2500 443.2000 ;
      RECT 432.9500 440.2000 438.1000 443.2000 ;
      RECT 424.8000 440.2000 429.9500 443.2000 ;
      RECT 416.6500 440.2000 421.8000 443.2000 ;
      RECT 396.5000 440.2000 413.6500 443.2000 ;
      RECT 346.5000 440.2000 393.5000 443.2000 ;
      RECT 326.4650 440.2000 343.5000 443.2000 ;
      RECT 317.9500 440.2000 323.4650 443.2000 ;
      RECT 309.4350 440.2000 314.9500 443.2000 ;
      RECT 300.9200 440.2000 306.4350 443.2000 ;
      RECT 292.4050 440.2000 297.9200 443.2000 ;
      RECT 283.8900 440.2000 289.4050 443.2000 ;
      RECT 275.3750 440.2000 280.8900 443.2000 ;
      RECT 266.8600 440.2000 272.3750 443.2000 ;
      RECT 258.3450 440.2000 263.8600 443.2000 ;
      RECT 249.8300 440.2000 255.3450 443.2000 ;
      RECT 241.3150 440.2000 246.8300 443.2000 ;
      RECT 232.8000 440.2000 238.3150 443.2000 ;
      RECT 224.2850 440.2000 229.8000 443.2000 ;
      RECT 215.7700 440.2000 221.2850 443.2000 ;
      RECT 207.2550 440.2000 212.7700 443.2000 ;
      RECT 198.7400 440.2000 204.2550 443.2000 ;
      RECT 190.2250 440.2000 195.7400 443.2000 ;
      RECT 181.7100 440.2000 187.2250 443.2000 ;
      RECT 173.1950 440.2000 178.7100 443.2000 ;
      RECT 164.6800 440.2000 170.1950 443.2000 ;
      RECT 156.1650 440.2000 161.6800 443.2000 ;
      RECT 147.6500 440.2000 153.1650 443.2000 ;
      RECT 139.1350 440.2000 144.6500 443.2000 ;
      RECT 130.6200 440.2000 136.1350 443.2000 ;
      RECT 122.1050 440.2000 127.6200 443.2000 ;
      RECT 113.5900 440.2000 119.1050 443.2000 ;
      RECT 105.0750 440.2000 110.5900 443.2000 ;
      RECT 96.5600 440.2000 102.0750 443.2000 ;
      RECT 88.0450 440.2000 93.5600 443.2000 ;
      RECT 79.5300 440.2000 85.0450 443.2000 ;
      RECT 71.0150 440.2000 76.5300 443.2000 ;
      RECT 62.5000 440.2000 68.0150 443.2000 ;
      RECT 46.5000 440.2000 59.5000 443.2000 ;
      RECT 8.5000 440.2000 43.5000 443.2000 ;
      RECT 0.0000 440.2000 5.5000 443.2000 ;
      RECT 0.0000 438.7000 1120.0000 440.2000 ;
      RECT 1116.6000 438.2000 1120.0000 438.7000 ;
      RECT 0.0000 436.1050 1113.6000 438.7000 ;
      RECT 1118.5000 435.2000 1120.0000 438.2000 ;
      RECT 1114.5000 433.1050 1120.0000 435.2000 ;
      RECT 1076.5000 433.1050 1111.5000 436.1050 ;
      RECT 1060.5000 433.1050 1073.5000 436.1050 ;
      RECT 1052.3500 433.1050 1057.5000 436.1050 ;
      RECT 1044.2000 433.1050 1049.3500 436.1050 ;
      RECT 1036.0500 433.1050 1041.2000 436.1050 ;
      RECT 1027.9000 433.1050 1033.0500 436.1050 ;
      RECT 1019.7500 433.1050 1024.9000 436.1050 ;
      RECT 1011.6000 433.1050 1016.7500 436.1050 ;
      RECT 1003.4500 433.1050 1008.6000 436.1050 ;
      RECT 995.3000 433.1050 1000.4500 436.1050 ;
      RECT 987.1500 433.1050 992.3000 436.1050 ;
      RECT 979.0000 433.1050 984.1500 436.1050 ;
      RECT 970.8500 433.1050 976.0000 436.1050 ;
      RECT 962.7000 433.1050 967.8500 436.1050 ;
      RECT 954.5500 433.1050 959.7000 436.1050 ;
      RECT 946.4000 433.1050 951.5500 436.1050 ;
      RECT 938.2500 433.1050 943.4000 436.1050 ;
      RECT 930.1000 433.1050 935.2500 436.1050 ;
      RECT 921.9500 433.1050 927.1000 436.1050 ;
      RECT 913.8000 433.1050 918.9500 436.1050 ;
      RECT 905.6500 433.1050 910.8000 436.1050 ;
      RECT 897.5000 433.1050 902.6500 436.1050 ;
      RECT 889.3500 433.1050 894.5000 436.1050 ;
      RECT 881.2000 433.1050 886.3500 436.1050 ;
      RECT 873.0500 433.1050 878.2000 436.1050 ;
      RECT 864.9000 433.1050 870.0500 436.1050 ;
      RECT 856.7500 433.1050 861.9000 436.1050 ;
      RECT 848.6000 433.1050 853.7500 436.1050 ;
      RECT 840.4500 433.1050 845.6000 436.1050 ;
      RECT 832.3000 433.1050 837.4500 436.1050 ;
      RECT 824.1500 433.1050 829.3000 436.1050 ;
      RECT 816.0000 433.1050 821.1500 436.1050 ;
      RECT 807.8500 433.1050 813.0000 436.1050 ;
      RECT 799.7000 433.1050 804.8500 436.1050 ;
      RECT 791.5500 433.1050 796.7000 436.1050 ;
      RECT 783.4000 433.1050 788.5500 436.1050 ;
      RECT 775.2500 433.1050 780.4000 436.1050 ;
      RECT 767.1000 433.1050 772.2500 436.1050 ;
      RECT 758.9500 433.1050 764.1000 436.1050 ;
      RECT 750.8000 433.1050 755.9500 436.1050 ;
      RECT 742.6500 433.1050 747.8000 436.1050 ;
      RECT 734.5000 433.1050 739.6500 436.1050 ;
      RECT 726.3500 433.1050 731.5000 436.1050 ;
      RECT 718.2000 433.1050 723.3500 436.1050 ;
      RECT 710.0500 433.1050 715.2000 436.1050 ;
      RECT 701.9000 433.1050 707.0500 436.1050 ;
      RECT 693.7500 433.1050 698.9000 436.1050 ;
      RECT 685.6000 433.1050 690.7500 436.1050 ;
      RECT 677.4500 433.1050 682.6000 436.1050 ;
      RECT 669.3000 433.1050 674.4500 436.1050 ;
      RECT 661.1500 433.1050 666.3000 436.1050 ;
      RECT 653.0000 433.1050 658.1500 436.1050 ;
      RECT 644.8500 433.1050 650.0000 436.1050 ;
      RECT 636.7000 433.1050 641.8500 436.1050 ;
      RECT 628.5500 433.1050 633.7000 436.1050 ;
      RECT 620.4000 433.1050 625.5500 436.1050 ;
      RECT 612.2500 433.1050 617.4000 436.1050 ;
      RECT 604.1000 433.1050 609.2500 436.1050 ;
      RECT 595.9500 433.1050 601.1000 436.1050 ;
      RECT 587.8000 433.1050 592.9500 436.1050 ;
      RECT 579.6500 433.1050 584.8000 436.1050 ;
      RECT 571.5000 433.1050 576.6500 436.1050 ;
      RECT 563.3500 433.1050 568.5000 436.1050 ;
      RECT 555.2000 433.1050 560.3500 436.1050 ;
      RECT 547.0500 433.1050 552.2000 436.1050 ;
      RECT 538.9000 433.1050 544.0500 436.1050 ;
      RECT 530.7500 433.1050 535.9000 436.1050 ;
      RECT 522.6000 433.1050 527.7500 436.1050 ;
      RECT 514.4500 433.1050 519.6000 436.1050 ;
      RECT 506.3000 433.1050 511.4500 436.1050 ;
      RECT 498.1500 433.1050 503.3000 436.1050 ;
      RECT 490.0000 433.1050 495.1500 436.1050 ;
      RECT 481.8500 433.1050 487.0000 436.1050 ;
      RECT 473.7000 433.1050 478.8500 436.1050 ;
      RECT 465.5500 433.1050 470.7000 436.1050 ;
      RECT 457.4000 433.1050 462.5500 436.1050 ;
      RECT 449.2500 433.1050 454.4000 436.1050 ;
      RECT 441.1000 433.1050 446.2500 436.1050 ;
      RECT 432.9500 433.1050 438.1000 436.1050 ;
      RECT 424.8000 433.1050 429.9500 436.1050 ;
      RECT 416.6500 433.1050 421.8000 436.1050 ;
      RECT 396.5000 433.1050 413.6500 436.1050 ;
      RECT 346.5000 433.1050 393.5000 436.1050 ;
      RECT 326.4650 433.1050 343.5000 436.1050 ;
      RECT 317.9500 433.1050 323.4650 436.1050 ;
      RECT 309.4350 433.1050 314.9500 436.1050 ;
      RECT 300.9200 433.1050 306.4350 436.1050 ;
      RECT 292.4050 433.1050 297.9200 436.1050 ;
      RECT 283.8900 433.1050 289.4050 436.1050 ;
      RECT 275.3750 433.1050 280.8900 436.1050 ;
      RECT 266.8600 433.1050 272.3750 436.1050 ;
      RECT 258.3450 433.1050 263.8600 436.1050 ;
      RECT 249.8300 433.1050 255.3450 436.1050 ;
      RECT 241.3150 433.1050 246.8300 436.1050 ;
      RECT 232.8000 433.1050 238.3150 436.1050 ;
      RECT 224.2850 433.1050 229.8000 436.1050 ;
      RECT 215.7700 433.1050 221.2850 436.1050 ;
      RECT 207.2550 433.1050 212.7700 436.1050 ;
      RECT 198.7400 433.1050 204.2550 436.1050 ;
      RECT 190.2250 433.1050 195.7400 436.1050 ;
      RECT 181.7100 433.1050 187.2250 436.1050 ;
      RECT 173.1950 433.1050 178.7100 436.1050 ;
      RECT 164.6800 433.1050 170.1950 436.1050 ;
      RECT 156.1650 433.1050 161.6800 436.1050 ;
      RECT 147.6500 433.1050 153.1650 436.1050 ;
      RECT 139.1350 433.1050 144.6500 436.1050 ;
      RECT 130.6200 433.1050 136.1350 436.1050 ;
      RECT 122.1050 433.1050 127.6200 436.1050 ;
      RECT 113.5900 433.1050 119.1050 436.1050 ;
      RECT 105.0750 433.1050 110.5900 436.1050 ;
      RECT 96.5600 433.1050 102.0750 436.1050 ;
      RECT 88.0450 433.1050 93.5600 436.1050 ;
      RECT 79.5300 433.1050 85.0450 436.1050 ;
      RECT 71.0150 433.1050 76.5300 436.1050 ;
      RECT 62.5000 433.1050 68.0150 436.1050 ;
      RECT 46.5000 433.1050 59.5000 436.1050 ;
      RECT 8.5000 433.1050 43.5000 436.1050 ;
      RECT 0.0000 433.1050 5.5000 436.1050 ;
      RECT 0.0000 431.7000 1120.0000 433.1050 ;
      RECT 1116.6000 431.1050 1120.0000 431.7000 ;
      RECT 0.0000 429.0100 1113.6000 431.7000 ;
      RECT 1118.5000 428.1050 1120.0000 431.1050 ;
      RECT 1114.5000 426.0100 1120.0000 428.1050 ;
      RECT 1076.5000 426.0100 1111.5000 429.0100 ;
      RECT 1060.5000 426.0100 1073.5000 429.0100 ;
      RECT 1052.3500 426.0100 1057.5000 429.0100 ;
      RECT 1044.2000 426.0100 1049.3500 429.0100 ;
      RECT 1036.0500 426.0100 1041.2000 429.0100 ;
      RECT 1027.9000 426.0100 1033.0500 429.0100 ;
      RECT 1019.7500 426.0100 1024.9000 429.0100 ;
      RECT 1011.6000 426.0100 1016.7500 429.0100 ;
      RECT 1003.4500 426.0100 1008.6000 429.0100 ;
      RECT 995.3000 426.0100 1000.4500 429.0100 ;
      RECT 987.1500 426.0100 992.3000 429.0100 ;
      RECT 979.0000 426.0100 984.1500 429.0100 ;
      RECT 970.8500 426.0100 976.0000 429.0100 ;
      RECT 962.7000 426.0100 967.8500 429.0100 ;
      RECT 954.5500 426.0100 959.7000 429.0100 ;
      RECT 946.4000 426.0100 951.5500 429.0100 ;
      RECT 938.2500 426.0100 943.4000 429.0100 ;
      RECT 930.1000 426.0100 935.2500 429.0100 ;
      RECT 921.9500 426.0100 927.1000 429.0100 ;
      RECT 913.8000 426.0100 918.9500 429.0100 ;
      RECT 905.6500 426.0100 910.8000 429.0100 ;
      RECT 897.5000 426.0100 902.6500 429.0100 ;
      RECT 889.3500 426.0100 894.5000 429.0100 ;
      RECT 881.2000 426.0100 886.3500 429.0100 ;
      RECT 873.0500 426.0100 878.2000 429.0100 ;
      RECT 864.9000 426.0100 870.0500 429.0100 ;
      RECT 856.7500 426.0100 861.9000 429.0100 ;
      RECT 848.6000 426.0100 853.7500 429.0100 ;
      RECT 840.4500 426.0100 845.6000 429.0100 ;
      RECT 832.3000 426.0100 837.4500 429.0100 ;
      RECT 824.1500 426.0100 829.3000 429.0100 ;
      RECT 816.0000 426.0100 821.1500 429.0100 ;
      RECT 807.8500 426.0100 813.0000 429.0100 ;
      RECT 799.7000 426.0100 804.8500 429.0100 ;
      RECT 791.5500 426.0100 796.7000 429.0100 ;
      RECT 783.4000 426.0100 788.5500 429.0100 ;
      RECT 775.2500 426.0100 780.4000 429.0100 ;
      RECT 767.1000 426.0100 772.2500 429.0100 ;
      RECT 758.9500 426.0100 764.1000 429.0100 ;
      RECT 750.8000 426.0100 755.9500 429.0100 ;
      RECT 742.6500 426.0100 747.8000 429.0100 ;
      RECT 734.5000 426.0100 739.6500 429.0100 ;
      RECT 726.3500 426.0100 731.5000 429.0100 ;
      RECT 718.2000 426.0100 723.3500 429.0100 ;
      RECT 710.0500 426.0100 715.2000 429.0100 ;
      RECT 701.9000 426.0100 707.0500 429.0100 ;
      RECT 693.7500 426.0100 698.9000 429.0100 ;
      RECT 685.6000 426.0100 690.7500 429.0100 ;
      RECT 677.4500 426.0100 682.6000 429.0100 ;
      RECT 669.3000 426.0100 674.4500 429.0100 ;
      RECT 661.1500 426.0100 666.3000 429.0100 ;
      RECT 653.0000 426.0100 658.1500 429.0100 ;
      RECT 644.8500 426.0100 650.0000 429.0100 ;
      RECT 636.7000 426.0100 641.8500 429.0100 ;
      RECT 628.5500 426.0100 633.7000 429.0100 ;
      RECT 620.4000 426.0100 625.5500 429.0100 ;
      RECT 612.2500 426.0100 617.4000 429.0100 ;
      RECT 604.1000 426.0100 609.2500 429.0100 ;
      RECT 595.9500 426.0100 601.1000 429.0100 ;
      RECT 587.8000 426.0100 592.9500 429.0100 ;
      RECT 579.6500 426.0100 584.8000 429.0100 ;
      RECT 571.5000 426.0100 576.6500 429.0100 ;
      RECT 563.3500 426.0100 568.5000 429.0100 ;
      RECT 555.2000 426.0100 560.3500 429.0100 ;
      RECT 547.0500 426.0100 552.2000 429.0100 ;
      RECT 538.9000 426.0100 544.0500 429.0100 ;
      RECT 530.7500 426.0100 535.9000 429.0100 ;
      RECT 522.6000 426.0100 527.7500 429.0100 ;
      RECT 514.4500 426.0100 519.6000 429.0100 ;
      RECT 506.3000 426.0100 511.4500 429.0100 ;
      RECT 498.1500 426.0100 503.3000 429.0100 ;
      RECT 490.0000 426.0100 495.1500 429.0100 ;
      RECT 481.8500 426.0100 487.0000 429.0100 ;
      RECT 473.7000 426.0100 478.8500 429.0100 ;
      RECT 465.5500 426.0100 470.7000 429.0100 ;
      RECT 457.4000 426.0100 462.5500 429.0100 ;
      RECT 449.2500 426.0100 454.4000 429.0100 ;
      RECT 441.1000 426.0100 446.2500 429.0100 ;
      RECT 432.9500 426.0100 438.1000 429.0100 ;
      RECT 424.8000 426.0100 429.9500 429.0100 ;
      RECT 416.6500 426.0100 421.8000 429.0100 ;
      RECT 396.5000 426.0100 413.6500 429.0100 ;
      RECT 346.5000 426.0100 393.5000 429.0100 ;
      RECT 326.4650 426.0100 343.5000 429.0100 ;
      RECT 317.9500 426.0100 323.4650 429.0100 ;
      RECT 309.4350 426.0100 314.9500 429.0100 ;
      RECT 300.9200 426.0100 306.4350 429.0100 ;
      RECT 292.4050 426.0100 297.9200 429.0100 ;
      RECT 283.8900 426.0100 289.4050 429.0100 ;
      RECT 275.3750 426.0100 280.8900 429.0100 ;
      RECT 266.8600 426.0100 272.3750 429.0100 ;
      RECT 258.3450 426.0100 263.8600 429.0100 ;
      RECT 249.8300 426.0100 255.3450 429.0100 ;
      RECT 241.3150 426.0100 246.8300 429.0100 ;
      RECT 232.8000 426.0100 238.3150 429.0100 ;
      RECT 224.2850 426.0100 229.8000 429.0100 ;
      RECT 215.7700 426.0100 221.2850 429.0100 ;
      RECT 207.2550 426.0100 212.7700 429.0100 ;
      RECT 198.7400 426.0100 204.2550 429.0100 ;
      RECT 190.2250 426.0100 195.7400 429.0100 ;
      RECT 181.7100 426.0100 187.2250 429.0100 ;
      RECT 173.1950 426.0100 178.7100 429.0100 ;
      RECT 164.6800 426.0100 170.1950 429.0100 ;
      RECT 156.1650 426.0100 161.6800 429.0100 ;
      RECT 147.6500 426.0100 153.1650 429.0100 ;
      RECT 139.1350 426.0100 144.6500 429.0100 ;
      RECT 130.6200 426.0100 136.1350 429.0100 ;
      RECT 122.1050 426.0100 127.6200 429.0100 ;
      RECT 113.5900 426.0100 119.1050 429.0100 ;
      RECT 105.0750 426.0100 110.5900 429.0100 ;
      RECT 96.5600 426.0100 102.0750 429.0100 ;
      RECT 88.0450 426.0100 93.5600 429.0100 ;
      RECT 79.5300 426.0100 85.0450 429.0100 ;
      RECT 71.0150 426.0100 76.5300 429.0100 ;
      RECT 62.5000 426.0100 68.0150 429.0100 ;
      RECT 46.5000 426.0100 59.5000 429.0100 ;
      RECT 8.5000 426.0100 43.5000 429.0100 ;
      RECT 0.0000 426.0100 5.5000 429.0100 ;
      RECT 0.0000 424.5000 1120.0000 426.0100 ;
      RECT 1116.6000 424.0100 1120.0000 424.5000 ;
      RECT 0.0000 421.9150 1113.6000 424.5000 ;
      RECT 1118.5000 421.0100 1120.0000 424.0100 ;
      RECT 1114.5000 418.9150 1120.0000 421.0100 ;
      RECT 1076.5000 418.9150 1111.5000 421.9150 ;
      RECT 1060.5000 418.9150 1073.5000 421.9150 ;
      RECT 1052.3500 418.9150 1057.5000 421.9150 ;
      RECT 1044.2000 418.9150 1049.3500 421.9150 ;
      RECT 1036.0500 418.9150 1041.2000 421.9150 ;
      RECT 1027.9000 418.9150 1033.0500 421.9150 ;
      RECT 1019.7500 418.9150 1024.9000 421.9150 ;
      RECT 1011.6000 418.9150 1016.7500 421.9150 ;
      RECT 1003.4500 418.9150 1008.6000 421.9150 ;
      RECT 995.3000 418.9150 1000.4500 421.9150 ;
      RECT 987.1500 418.9150 992.3000 421.9150 ;
      RECT 979.0000 418.9150 984.1500 421.9150 ;
      RECT 970.8500 418.9150 976.0000 421.9150 ;
      RECT 962.7000 418.9150 967.8500 421.9150 ;
      RECT 954.5500 418.9150 959.7000 421.9150 ;
      RECT 946.4000 418.9150 951.5500 421.9150 ;
      RECT 938.2500 418.9150 943.4000 421.9150 ;
      RECT 930.1000 418.9150 935.2500 421.9150 ;
      RECT 921.9500 418.9150 927.1000 421.9150 ;
      RECT 913.8000 418.9150 918.9500 421.9150 ;
      RECT 905.6500 418.9150 910.8000 421.9150 ;
      RECT 897.5000 418.9150 902.6500 421.9150 ;
      RECT 889.3500 418.9150 894.5000 421.9150 ;
      RECT 881.2000 418.9150 886.3500 421.9150 ;
      RECT 873.0500 418.9150 878.2000 421.9150 ;
      RECT 864.9000 418.9150 870.0500 421.9150 ;
      RECT 856.7500 418.9150 861.9000 421.9150 ;
      RECT 848.6000 418.9150 853.7500 421.9150 ;
      RECT 840.4500 418.9150 845.6000 421.9150 ;
      RECT 832.3000 418.9150 837.4500 421.9150 ;
      RECT 824.1500 418.9150 829.3000 421.9150 ;
      RECT 816.0000 418.9150 821.1500 421.9150 ;
      RECT 807.8500 418.9150 813.0000 421.9150 ;
      RECT 799.7000 418.9150 804.8500 421.9150 ;
      RECT 791.5500 418.9150 796.7000 421.9150 ;
      RECT 783.4000 418.9150 788.5500 421.9150 ;
      RECT 775.2500 418.9150 780.4000 421.9150 ;
      RECT 767.1000 418.9150 772.2500 421.9150 ;
      RECT 758.9500 418.9150 764.1000 421.9150 ;
      RECT 750.8000 418.9150 755.9500 421.9150 ;
      RECT 742.6500 418.9150 747.8000 421.9150 ;
      RECT 734.5000 418.9150 739.6500 421.9150 ;
      RECT 726.3500 418.9150 731.5000 421.9150 ;
      RECT 718.2000 418.9150 723.3500 421.9150 ;
      RECT 710.0500 418.9150 715.2000 421.9150 ;
      RECT 701.9000 418.9150 707.0500 421.9150 ;
      RECT 693.7500 418.9150 698.9000 421.9150 ;
      RECT 685.6000 418.9150 690.7500 421.9150 ;
      RECT 677.4500 418.9150 682.6000 421.9150 ;
      RECT 669.3000 418.9150 674.4500 421.9150 ;
      RECT 661.1500 418.9150 666.3000 421.9150 ;
      RECT 653.0000 418.9150 658.1500 421.9150 ;
      RECT 644.8500 418.9150 650.0000 421.9150 ;
      RECT 636.7000 418.9150 641.8500 421.9150 ;
      RECT 628.5500 418.9150 633.7000 421.9150 ;
      RECT 620.4000 418.9150 625.5500 421.9150 ;
      RECT 612.2500 418.9150 617.4000 421.9150 ;
      RECT 604.1000 418.9150 609.2500 421.9150 ;
      RECT 595.9500 418.9150 601.1000 421.9150 ;
      RECT 587.8000 418.9150 592.9500 421.9150 ;
      RECT 579.6500 418.9150 584.8000 421.9150 ;
      RECT 571.5000 418.9150 576.6500 421.9150 ;
      RECT 563.3500 418.9150 568.5000 421.9150 ;
      RECT 555.2000 418.9150 560.3500 421.9150 ;
      RECT 547.0500 418.9150 552.2000 421.9150 ;
      RECT 538.9000 418.9150 544.0500 421.9150 ;
      RECT 530.7500 418.9150 535.9000 421.9150 ;
      RECT 522.6000 418.9150 527.7500 421.9150 ;
      RECT 514.4500 418.9150 519.6000 421.9150 ;
      RECT 506.3000 418.9150 511.4500 421.9150 ;
      RECT 498.1500 418.9150 503.3000 421.9150 ;
      RECT 490.0000 418.9150 495.1500 421.9150 ;
      RECT 481.8500 418.9150 487.0000 421.9150 ;
      RECT 473.7000 418.9150 478.8500 421.9150 ;
      RECT 465.5500 418.9150 470.7000 421.9150 ;
      RECT 457.4000 418.9150 462.5500 421.9150 ;
      RECT 449.2500 418.9150 454.4000 421.9150 ;
      RECT 441.1000 418.9150 446.2500 421.9150 ;
      RECT 432.9500 418.9150 438.1000 421.9150 ;
      RECT 424.8000 418.9150 429.9500 421.9150 ;
      RECT 416.6500 418.9150 421.8000 421.9150 ;
      RECT 396.5000 418.9150 413.6500 421.9150 ;
      RECT 346.5000 418.9150 393.5000 421.9150 ;
      RECT 326.4650 418.9150 343.5000 421.9150 ;
      RECT 317.9500 418.9150 323.4650 421.9150 ;
      RECT 309.4350 418.9150 314.9500 421.9150 ;
      RECT 300.9200 418.9150 306.4350 421.9150 ;
      RECT 292.4050 418.9150 297.9200 421.9150 ;
      RECT 283.8900 418.9150 289.4050 421.9150 ;
      RECT 275.3750 418.9150 280.8900 421.9150 ;
      RECT 266.8600 418.9150 272.3750 421.9150 ;
      RECT 258.3450 418.9150 263.8600 421.9150 ;
      RECT 249.8300 418.9150 255.3450 421.9150 ;
      RECT 241.3150 418.9150 246.8300 421.9150 ;
      RECT 232.8000 418.9150 238.3150 421.9150 ;
      RECT 224.2850 418.9150 229.8000 421.9150 ;
      RECT 215.7700 418.9150 221.2850 421.9150 ;
      RECT 207.2550 418.9150 212.7700 421.9150 ;
      RECT 198.7400 418.9150 204.2550 421.9150 ;
      RECT 190.2250 418.9150 195.7400 421.9150 ;
      RECT 181.7100 418.9150 187.2250 421.9150 ;
      RECT 173.1950 418.9150 178.7100 421.9150 ;
      RECT 164.6800 418.9150 170.1950 421.9150 ;
      RECT 156.1650 418.9150 161.6800 421.9150 ;
      RECT 147.6500 418.9150 153.1650 421.9150 ;
      RECT 139.1350 418.9150 144.6500 421.9150 ;
      RECT 130.6200 418.9150 136.1350 421.9150 ;
      RECT 122.1050 418.9150 127.6200 421.9150 ;
      RECT 113.5900 418.9150 119.1050 421.9150 ;
      RECT 105.0750 418.9150 110.5900 421.9150 ;
      RECT 96.5600 418.9150 102.0750 421.9150 ;
      RECT 88.0450 418.9150 93.5600 421.9150 ;
      RECT 79.5300 418.9150 85.0450 421.9150 ;
      RECT 71.0150 418.9150 76.5300 421.9150 ;
      RECT 62.5000 418.9150 68.0150 421.9150 ;
      RECT 46.5000 418.9150 59.5000 421.9150 ;
      RECT 8.5000 418.9150 43.5000 421.9150 ;
      RECT 0.0000 418.9150 5.5000 421.9150 ;
      RECT 0.0000 417.5000 1120.0000 418.9150 ;
      RECT 1116.6000 416.9150 1120.0000 417.5000 ;
      RECT 0.0000 414.8200 1113.6000 417.5000 ;
      RECT 1118.5000 413.9150 1120.0000 416.9150 ;
      RECT 1114.5000 411.8200 1120.0000 413.9150 ;
      RECT 1076.5000 411.8200 1111.5000 414.8200 ;
      RECT 1060.5000 411.8200 1073.5000 414.8200 ;
      RECT 1052.3500 411.8200 1057.5000 414.8200 ;
      RECT 1044.2000 411.8200 1049.3500 414.8200 ;
      RECT 1036.0500 411.8200 1041.2000 414.8200 ;
      RECT 1027.9000 411.8200 1033.0500 414.8200 ;
      RECT 1019.7500 411.8200 1024.9000 414.8200 ;
      RECT 1011.6000 411.8200 1016.7500 414.8200 ;
      RECT 1003.4500 411.8200 1008.6000 414.8200 ;
      RECT 995.3000 411.8200 1000.4500 414.8200 ;
      RECT 987.1500 411.8200 992.3000 414.8200 ;
      RECT 979.0000 411.8200 984.1500 414.8200 ;
      RECT 970.8500 411.8200 976.0000 414.8200 ;
      RECT 962.7000 411.8200 967.8500 414.8200 ;
      RECT 954.5500 411.8200 959.7000 414.8200 ;
      RECT 946.4000 411.8200 951.5500 414.8200 ;
      RECT 938.2500 411.8200 943.4000 414.8200 ;
      RECT 930.1000 411.8200 935.2500 414.8200 ;
      RECT 921.9500 411.8200 927.1000 414.8200 ;
      RECT 913.8000 411.8200 918.9500 414.8200 ;
      RECT 905.6500 411.8200 910.8000 414.8200 ;
      RECT 897.5000 411.8200 902.6500 414.8200 ;
      RECT 889.3500 411.8200 894.5000 414.8200 ;
      RECT 881.2000 411.8200 886.3500 414.8200 ;
      RECT 873.0500 411.8200 878.2000 414.8200 ;
      RECT 864.9000 411.8200 870.0500 414.8200 ;
      RECT 856.7500 411.8200 861.9000 414.8200 ;
      RECT 848.6000 411.8200 853.7500 414.8200 ;
      RECT 840.4500 411.8200 845.6000 414.8200 ;
      RECT 832.3000 411.8200 837.4500 414.8200 ;
      RECT 824.1500 411.8200 829.3000 414.8200 ;
      RECT 816.0000 411.8200 821.1500 414.8200 ;
      RECT 807.8500 411.8200 813.0000 414.8200 ;
      RECT 799.7000 411.8200 804.8500 414.8200 ;
      RECT 791.5500 411.8200 796.7000 414.8200 ;
      RECT 783.4000 411.8200 788.5500 414.8200 ;
      RECT 775.2500 411.8200 780.4000 414.8200 ;
      RECT 767.1000 411.8200 772.2500 414.8200 ;
      RECT 758.9500 411.8200 764.1000 414.8200 ;
      RECT 750.8000 411.8200 755.9500 414.8200 ;
      RECT 742.6500 411.8200 747.8000 414.8200 ;
      RECT 734.5000 411.8200 739.6500 414.8200 ;
      RECT 726.3500 411.8200 731.5000 414.8200 ;
      RECT 718.2000 411.8200 723.3500 414.8200 ;
      RECT 710.0500 411.8200 715.2000 414.8200 ;
      RECT 701.9000 411.8200 707.0500 414.8200 ;
      RECT 693.7500 411.8200 698.9000 414.8200 ;
      RECT 685.6000 411.8200 690.7500 414.8200 ;
      RECT 677.4500 411.8200 682.6000 414.8200 ;
      RECT 669.3000 411.8200 674.4500 414.8200 ;
      RECT 661.1500 411.8200 666.3000 414.8200 ;
      RECT 653.0000 411.8200 658.1500 414.8200 ;
      RECT 644.8500 411.8200 650.0000 414.8200 ;
      RECT 636.7000 411.8200 641.8500 414.8200 ;
      RECT 628.5500 411.8200 633.7000 414.8200 ;
      RECT 620.4000 411.8200 625.5500 414.8200 ;
      RECT 612.2500 411.8200 617.4000 414.8200 ;
      RECT 604.1000 411.8200 609.2500 414.8200 ;
      RECT 595.9500 411.8200 601.1000 414.8200 ;
      RECT 587.8000 411.8200 592.9500 414.8200 ;
      RECT 579.6500 411.8200 584.8000 414.8200 ;
      RECT 571.5000 411.8200 576.6500 414.8200 ;
      RECT 563.3500 411.8200 568.5000 414.8200 ;
      RECT 555.2000 411.8200 560.3500 414.8200 ;
      RECT 547.0500 411.8200 552.2000 414.8200 ;
      RECT 538.9000 411.8200 544.0500 414.8200 ;
      RECT 530.7500 411.8200 535.9000 414.8200 ;
      RECT 522.6000 411.8200 527.7500 414.8200 ;
      RECT 514.4500 411.8200 519.6000 414.8200 ;
      RECT 506.3000 411.8200 511.4500 414.8200 ;
      RECT 498.1500 411.8200 503.3000 414.8200 ;
      RECT 490.0000 411.8200 495.1500 414.8200 ;
      RECT 481.8500 411.8200 487.0000 414.8200 ;
      RECT 473.7000 411.8200 478.8500 414.8200 ;
      RECT 465.5500 411.8200 470.7000 414.8200 ;
      RECT 457.4000 411.8200 462.5500 414.8200 ;
      RECT 449.2500 411.8200 454.4000 414.8200 ;
      RECT 441.1000 411.8200 446.2500 414.8200 ;
      RECT 432.9500 411.8200 438.1000 414.8200 ;
      RECT 424.8000 411.8200 429.9500 414.8200 ;
      RECT 416.6500 411.8200 421.8000 414.8200 ;
      RECT 396.5000 411.8200 413.6500 414.8200 ;
      RECT 346.5000 411.8200 393.5000 414.8200 ;
      RECT 326.4650 411.8200 343.5000 414.8200 ;
      RECT 317.9500 411.8200 323.4650 414.8200 ;
      RECT 309.4350 411.8200 314.9500 414.8200 ;
      RECT 300.9200 411.8200 306.4350 414.8200 ;
      RECT 292.4050 411.8200 297.9200 414.8200 ;
      RECT 283.8900 411.8200 289.4050 414.8200 ;
      RECT 275.3750 411.8200 280.8900 414.8200 ;
      RECT 266.8600 411.8200 272.3750 414.8200 ;
      RECT 258.3450 411.8200 263.8600 414.8200 ;
      RECT 249.8300 411.8200 255.3450 414.8200 ;
      RECT 241.3150 411.8200 246.8300 414.8200 ;
      RECT 232.8000 411.8200 238.3150 414.8200 ;
      RECT 224.2850 411.8200 229.8000 414.8200 ;
      RECT 215.7700 411.8200 221.2850 414.8200 ;
      RECT 207.2550 411.8200 212.7700 414.8200 ;
      RECT 198.7400 411.8200 204.2550 414.8200 ;
      RECT 190.2250 411.8200 195.7400 414.8200 ;
      RECT 181.7100 411.8200 187.2250 414.8200 ;
      RECT 173.1950 411.8200 178.7100 414.8200 ;
      RECT 164.6800 411.8200 170.1950 414.8200 ;
      RECT 156.1650 411.8200 161.6800 414.8200 ;
      RECT 147.6500 411.8200 153.1650 414.8200 ;
      RECT 139.1350 411.8200 144.6500 414.8200 ;
      RECT 130.6200 411.8200 136.1350 414.8200 ;
      RECT 122.1050 411.8200 127.6200 414.8200 ;
      RECT 113.5900 411.8200 119.1050 414.8200 ;
      RECT 105.0750 411.8200 110.5900 414.8200 ;
      RECT 96.5600 411.8200 102.0750 414.8200 ;
      RECT 88.0450 411.8200 93.5600 414.8200 ;
      RECT 79.5300 411.8200 85.0450 414.8200 ;
      RECT 71.0150 411.8200 76.5300 414.8200 ;
      RECT 62.5000 411.8200 68.0150 414.8200 ;
      RECT 46.5000 411.8200 59.5000 414.8200 ;
      RECT 8.5000 411.8200 43.5000 414.8200 ;
      RECT 0.0000 411.8200 5.5000 414.8200 ;
      RECT 0.0000 410.3000 1120.0000 411.8200 ;
      RECT 1116.6000 409.8200 1120.0000 410.3000 ;
      RECT 0.0000 407.7250 1113.6000 410.3000 ;
      RECT 1118.5000 406.8200 1120.0000 409.8200 ;
      RECT 1114.5000 404.7250 1120.0000 406.8200 ;
      RECT 1076.5000 404.7250 1111.5000 407.7250 ;
      RECT 1060.5000 404.7250 1073.5000 407.7250 ;
      RECT 1052.3500 404.7250 1057.5000 407.7250 ;
      RECT 1044.2000 404.7250 1049.3500 407.7250 ;
      RECT 1036.0500 404.7250 1041.2000 407.7250 ;
      RECT 1027.9000 404.7250 1033.0500 407.7250 ;
      RECT 1019.7500 404.7250 1024.9000 407.7250 ;
      RECT 1011.6000 404.7250 1016.7500 407.7250 ;
      RECT 1003.4500 404.7250 1008.6000 407.7250 ;
      RECT 995.3000 404.7250 1000.4500 407.7250 ;
      RECT 987.1500 404.7250 992.3000 407.7250 ;
      RECT 979.0000 404.7250 984.1500 407.7250 ;
      RECT 970.8500 404.7250 976.0000 407.7250 ;
      RECT 962.7000 404.7250 967.8500 407.7250 ;
      RECT 954.5500 404.7250 959.7000 407.7250 ;
      RECT 946.4000 404.7250 951.5500 407.7250 ;
      RECT 938.2500 404.7250 943.4000 407.7250 ;
      RECT 930.1000 404.7250 935.2500 407.7250 ;
      RECT 921.9500 404.7250 927.1000 407.7250 ;
      RECT 913.8000 404.7250 918.9500 407.7250 ;
      RECT 905.6500 404.7250 910.8000 407.7250 ;
      RECT 897.5000 404.7250 902.6500 407.7250 ;
      RECT 889.3500 404.7250 894.5000 407.7250 ;
      RECT 881.2000 404.7250 886.3500 407.7250 ;
      RECT 873.0500 404.7250 878.2000 407.7250 ;
      RECT 864.9000 404.7250 870.0500 407.7250 ;
      RECT 856.7500 404.7250 861.9000 407.7250 ;
      RECT 848.6000 404.7250 853.7500 407.7250 ;
      RECT 840.4500 404.7250 845.6000 407.7250 ;
      RECT 832.3000 404.7250 837.4500 407.7250 ;
      RECT 824.1500 404.7250 829.3000 407.7250 ;
      RECT 816.0000 404.7250 821.1500 407.7250 ;
      RECT 807.8500 404.7250 813.0000 407.7250 ;
      RECT 799.7000 404.7250 804.8500 407.7250 ;
      RECT 791.5500 404.7250 796.7000 407.7250 ;
      RECT 783.4000 404.7250 788.5500 407.7250 ;
      RECT 775.2500 404.7250 780.4000 407.7250 ;
      RECT 767.1000 404.7250 772.2500 407.7250 ;
      RECT 758.9500 404.7250 764.1000 407.7250 ;
      RECT 750.8000 404.7250 755.9500 407.7250 ;
      RECT 742.6500 404.7250 747.8000 407.7250 ;
      RECT 734.5000 404.7250 739.6500 407.7250 ;
      RECT 726.3500 404.7250 731.5000 407.7250 ;
      RECT 718.2000 404.7250 723.3500 407.7250 ;
      RECT 710.0500 404.7250 715.2000 407.7250 ;
      RECT 701.9000 404.7250 707.0500 407.7250 ;
      RECT 693.7500 404.7250 698.9000 407.7250 ;
      RECT 685.6000 404.7250 690.7500 407.7250 ;
      RECT 677.4500 404.7250 682.6000 407.7250 ;
      RECT 669.3000 404.7250 674.4500 407.7250 ;
      RECT 661.1500 404.7250 666.3000 407.7250 ;
      RECT 653.0000 404.7250 658.1500 407.7250 ;
      RECT 644.8500 404.7250 650.0000 407.7250 ;
      RECT 636.7000 404.7250 641.8500 407.7250 ;
      RECT 628.5500 404.7250 633.7000 407.7250 ;
      RECT 620.4000 404.7250 625.5500 407.7250 ;
      RECT 612.2500 404.7250 617.4000 407.7250 ;
      RECT 604.1000 404.7250 609.2500 407.7250 ;
      RECT 595.9500 404.7250 601.1000 407.7250 ;
      RECT 587.8000 404.7250 592.9500 407.7250 ;
      RECT 579.6500 404.7250 584.8000 407.7250 ;
      RECT 571.5000 404.7250 576.6500 407.7250 ;
      RECT 563.3500 404.7250 568.5000 407.7250 ;
      RECT 555.2000 404.7250 560.3500 407.7250 ;
      RECT 547.0500 404.7250 552.2000 407.7250 ;
      RECT 538.9000 404.7250 544.0500 407.7250 ;
      RECT 530.7500 404.7250 535.9000 407.7250 ;
      RECT 522.6000 404.7250 527.7500 407.7250 ;
      RECT 514.4500 404.7250 519.6000 407.7250 ;
      RECT 506.3000 404.7250 511.4500 407.7250 ;
      RECT 498.1500 404.7250 503.3000 407.7250 ;
      RECT 490.0000 404.7250 495.1500 407.7250 ;
      RECT 481.8500 404.7250 487.0000 407.7250 ;
      RECT 473.7000 404.7250 478.8500 407.7250 ;
      RECT 465.5500 404.7250 470.7000 407.7250 ;
      RECT 457.4000 404.7250 462.5500 407.7250 ;
      RECT 449.2500 404.7250 454.4000 407.7250 ;
      RECT 441.1000 404.7250 446.2500 407.7250 ;
      RECT 432.9500 404.7250 438.1000 407.7250 ;
      RECT 424.8000 404.7250 429.9500 407.7250 ;
      RECT 416.6500 404.7250 421.8000 407.7250 ;
      RECT 396.5000 404.7250 413.6500 407.7250 ;
      RECT 346.5000 404.7250 393.5000 407.7250 ;
      RECT 46.5000 404.7250 343.5000 407.7250 ;
      RECT 8.5000 404.7250 43.5000 407.7250 ;
      RECT 0.0000 404.7250 5.5000 407.7250 ;
      RECT 0.0000 403.3000 1120.0000 404.7250 ;
      RECT 1116.6000 402.7250 1120.0000 403.3000 ;
      RECT 0.0000 400.6300 1113.6000 403.3000 ;
      RECT 1118.5000 399.7250 1120.0000 402.7250 ;
      RECT 1114.5000 397.6300 1120.0000 399.7250 ;
      RECT 1076.5000 397.6300 1111.5000 400.6300 ;
      RECT 1060.5000 397.6300 1073.5000 400.6300 ;
      RECT 1052.3500 397.6300 1057.5000 400.6300 ;
      RECT 1044.2000 397.6300 1049.3500 400.6300 ;
      RECT 1036.0500 397.6300 1041.2000 400.6300 ;
      RECT 1027.9000 397.6300 1033.0500 400.6300 ;
      RECT 1019.7500 397.6300 1024.9000 400.6300 ;
      RECT 1011.6000 397.6300 1016.7500 400.6300 ;
      RECT 1003.4500 397.6300 1008.6000 400.6300 ;
      RECT 995.3000 397.6300 1000.4500 400.6300 ;
      RECT 987.1500 397.6300 992.3000 400.6300 ;
      RECT 979.0000 397.6300 984.1500 400.6300 ;
      RECT 970.8500 397.6300 976.0000 400.6300 ;
      RECT 962.7000 397.6300 967.8500 400.6300 ;
      RECT 954.5500 397.6300 959.7000 400.6300 ;
      RECT 946.4000 397.6300 951.5500 400.6300 ;
      RECT 938.2500 397.6300 943.4000 400.6300 ;
      RECT 930.1000 397.6300 935.2500 400.6300 ;
      RECT 921.9500 397.6300 927.1000 400.6300 ;
      RECT 913.8000 397.6300 918.9500 400.6300 ;
      RECT 905.6500 397.6300 910.8000 400.6300 ;
      RECT 897.5000 397.6300 902.6500 400.6300 ;
      RECT 889.3500 397.6300 894.5000 400.6300 ;
      RECT 881.2000 397.6300 886.3500 400.6300 ;
      RECT 873.0500 397.6300 878.2000 400.6300 ;
      RECT 864.9000 397.6300 870.0500 400.6300 ;
      RECT 856.7500 397.6300 861.9000 400.6300 ;
      RECT 848.6000 397.6300 853.7500 400.6300 ;
      RECT 840.4500 397.6300 845.6000 400.6300 ;
      RECT 832.3000 397.6300 837.4500 400.6300 ;
      RECT 824.1500 397.6300 829.3000 400.6300 ;
      RECT 816.0000 397.6300 821.1500 400.6300 ;
      RECT 807.8500 397.6300 813.0000 400.6300 ;
      RECT 799.7000 397.6300 804.8500 400.6300 ;
      RECT 791.5500 397.6300 796.7000 400.6300 ;
      RECT 783.4000 397.6300 788.5500 400.6300 ;
      RECT 775.2500 397.6300 780.4000 400.6300 ;
      RECT 767.1000 397.6300 772.2500 400.6300 ;
      RECT 758.9500 397.6300 764.1000 400.6300 ;
      RECT 750.8000 397.6300 755.9500 400.6300 ;
      RECT 742.6500 397.6300 747.8000 400.6300 ;
      RECT 734.5000 397.6300 739.6500 400.6300 ;
      RECT 726.3500 397.6300 731.5000 400.6300 ;
      RECT 718.2000 397.6300 723.3500 400.6300 ;
      RECT 710.0500 397.6300 715.2000 400.6300 ;
      RECT 701.9000 397.6300 707.0500 400.6300 ;
      RECT 693.7500 397.6300 698.9000 400.6300 ;
      RECT 685.6000 397.6300 690.7500 400.6300 ;
      RECT 677.4500 397.6300 682.6000 400.6300 ;
      RECT 669.3000 397.6300 674.4500 400.6300 ;
      RECT 661.1500 397.6300 666.3000 400.6300 ;
      RECT 653.0000 397.6300 658.1500 400.6300 ;
      RECT 644.8500 397.6300 650.0000 400.6300 ;
      RECT 636.7000 397.6300 641.8500 400.6300 ;
      RECT 628.5500 397.6300 633.7000 400.6300 ;
      RECT 620.4000 397.6300 625.5500 400.6300 ;
      RECT 612.2500 397.6300 617.4000 400.6300 ;
      RECT 604.1000 397.6300 609.2500 400.6300 ;
      RECT 595.9500 397.6300 601.1000 400.6300 ;
      RECT 587.8000 397.6300 592.9500 400.6300 ;
      RECT 579.6500 397.6300 584.8000 400.6300 ;
      RECT 571.5000 397.6300 576.6500 400.6300 ;
      RECT 563.3500 397.6300 568.5000 400.6300 ;
      RECT 555.2000 397.6300 560.3500 400.6300 ;
      RECT 547.0500 397.6300 552.2000 400.6300 ;
      RECT 538.9000 397.6300 544.0500 400.6300 ;
      RECT 530.7500 397.6300 535.9000 400.6300 ;
      RECT 522.6000 397.6300 527.7500 400.6300 ;
      RECT 514.4500 397.6300 519.6000 400.6300 ;
      RECT 506.3000 397.6300 511.4500 400.6300 ;
      RECT 498.1500 397.6300 503.3000 400.6300 ;
      RECT 490.0000 397.6300 495.1500 400.6300 ;
      RECT 481.8500 397.6300 487.0000 400.6300 ;
      RECT 473.7000 397.6300 478.8500 400.6300 ;
      RECT 465.5500 397.6300 470.7000 400.6300 ;
      RECT 457.4000 397.6300 462.5500 400.6300 ;
      RECT 449.2500 397.6300 454.4000 400.6300 ;
      RECT 441.1000 397.6300 446.2500 400.6300 ;
      RECT 432.9500 397.6300 438.1000 400.6300 ;
      RECT 424.8000 397.6300 429.9500 400.6300 ;
      RECT 416.6500 397.6300 421.8000 400.6300 ;
      RECT 396.5000 397.6300 413.6500 400.6300 ;
      RECT 346.5000 397.6300 393.5000 400.6300 ;
      RECT 46.5000 397.6300 343.5000 400.6300 ;
      RECT 8.5000 397.6300 43.5000 400.6300 ;
      RECT 0.0000 397.6300 5.5000 400.6300 ;
      RECT 0.0000 396.3000 1120.0000 397.6300 ;
      RECT 1116.6000 395.6300 1120.0000 396.3000 ;
      RECT 0.0000 393.5350 1113.6000 396.3000 ;
      RECT 1118.5000 392.6300 1120.0000 395.6300 ;
      RECT 1114.5000 390.5350 1120.0000 392.6300 ;
      RECT 1076.5000 390.5350 1111.5000 393.5350 ;
      RECT 1060.5000 390.5350 1073.5000 393.5350 ;
      RECT 1052.3500 390.5350 1057.5000 393.5350 ;
      RECT 1044.2000 390.5350 1049.3500 393.5350 ;
      RECT 1036.0500 390.5350 1041.2000 393.5350 ;
      RECT 1027.9000 390.5350 1033.0500 393.5350 ;
      RECT 1019.7500 390.5350 1024.9000 393.5350 ;
      RECT 1011.6000 390.5350 1016.7500 393.5350 ;
      RECT 1003.4500 390.5350 1008.6000 393.5350 ;
      RECT 995.3000 390.5350 1000.4500 393.5350 ;
      RECT 987.1500 390.5350 992.3000 393.5350 ;
      RECT 979.0000 390.5350 984.1500 393.5350 ;
      RECT 970.8500 390.5350 976.0000 393.5350 ;
      RECT 962.7000 390.5350 967.8500 393.5350 ;
      RECT 954.5500 390.5350 959.7000 393.5350 ;
      RECT 946.4000 390.5350 951.5500 393.5350 ;
      RECT 938.2500 390.5350 943.4000 393.5350 ;
      RECT 930.1000 390.5350 935.2500 393.5350 ;
      RECT 921.9500 390.5350 927.1000 393.5350 ;
      RECT 913.8000 390.5350 918.9500 393.5350 ;
      RECT 905.6500 390.5350 910.8000 393.5350 ;
      RECT 897.5000 390.5350 902.6500 393.5350 ;
      RECT 889.3500 390.5350 894.5000 393.5350 ;
      RECT 881.2000 390.5350 886.3500 393.5350 ;
      RECT 873.0500 390.5350 878.2000 393.5350 ;
      RECT 864.9000 390.5350 870.0500 393.5350 ;
      RECT 856.7500 390.5350 861.9000 393.5350 ;
      RECT 848.6000 390.5350 853.7500 393.5350 ;
      RECT 840.4500 390.5350 845.6000 393.5350 ;
      RECT 832.3000 390.5350 837.4500 393.5350 ;
      RECT 824.1500 390.5350 829.3000 393.5350 ;
      RECT 816.0000 390.5350 821.1500 393.5350 ;
      RECT 807.8500 390.5350 813.0000 393.5350 ;
      RECT 799.7000 390.5350 804.8500 393.5350 ;
      RECT 791.5500 390.5350 796.7000 393.5350 ;
      RECT 783.4000 390.5350 788.5500 393.5350 ;
      RECT 775.2500 390.5350 780.4000 393.5350 ;
      RECT 767.1000 390.5350 772.2500 393.5350 ;
      RECT 758.9500 390.5350 764.1000 393.5350 ;
      RECT 750.8000 390.5350 755.9500 393.5350 ;
      RECT 742.6500 390.5350 747.8000 393.5350 ;
      RECT 734.5000 390.5350 739.6500 393.5350 ;
      RECT 726.3500 390.5350 731.5000 393.5350 ;
      RECT 718.2000 390.5350 723.3500 393.5350 ;
      RECT 710.0500 390.5350 715.2000 393.5350 ;
      RECT 701.9000 390.5350 707.0500 393.5350 ;
      RECT 693.7500 390.5350 698.9000 393.5350 ;
      RECT 685.6000 390.5350 690.7500 393.5350 ;
      RECT 677.4500 390.5350 682.6000 393.5350 ;
      RECT 669.3000 390.5350 674.4500 393.5350 ;
      RECT 661.1500 390.5350 666.3000 393.5350 ;
      RECT 653.0000 390.5350 658.1500 393.5350 ;
      RECT 644.8500 390.5350 650.0000 393.5350 ;
      RECT 636.7000 390.5350 641.8500 393.5350 ;
      RECT 628.5500 390.5350 633.7000 393.5350 ;
      RECT 620.4000 390.5350 625.5500 393.5350 ;
      RECT 612.2500 390.5350 617.4000 393.5350 ;
      RECT 604.1000 390.5350 609.2500 393.5350 ;
      RECT 595.9500 390.5350 601.1000 393.5350 ;
      RECT 587.8000 390.5350 592.9500 393.5350 ;
      RECT 579.6500 390.5350 584.8000 393.5350 ;
      RECT 571.5000 390.5350 576.6500 393.5350 ;
      RECT 563.3500 390.5350 568.5000 393.5350 ;
      RECT 555.2000 390.5350 560.3500 393.5350 ;
      RECT 547.0500 390.5350 552.2000 393.5350 ;
      RECT 538.9000 390.5350 544.0500 393.5350 ;
      RECT 530.7500 390.5350 535.9000 393.5350 ;
      RECT 522.6000 390.5350 527.7500 393.5350 ;
      RECT 514.4500 390.5350 519.6000 393.5350 ;
      RECT 506.3000 390.5350 511.4500 393.5350 ;
      RECT 498.1500 390.5350 503.3000 393.5350 ;
      RECT 490.0000 390.5350 495.1500 393.5350 ;
      RECT 481.8500 390.5350 487.0000 393.5350 ;
      RECT 473.7000 390.5350 478.8500 393.5350 ;
      RECT 465.5500 390.5350 470.7000 393.5350 ;
      RECT 457.4000 390.5350 462.5500 393.5350 ;
      RECT 449.2500 390.5350 454.4000 393.5350 ;
      RECT 441.1000 390.5350 446.2500 393.5350 ;
      RECT 432.9500 390.5350 438.1000 393.5350 ;
      RECT 424.8000 390.5350 429.9500 393.5350 ;
      RECT 416.6500 390.5350 421.8000 393.5350 ;
      RECT 396.5000 390.5350 413.6500 393.5350 ;
      RECT 8.5000 390.5350 393.5000 393.5350 ;
      RECT 0.0000 390.5350 5.5000 393.5350 ;
      RECT 0.0000 389.1000 1120.0000 390.5350 ;
      RECT 1116.6000 388.5350 1120.0000 389.1000 ;
      RECT 0.0000 386.4400 1113.6000 389.1000 ;
      RECT 1118.5000 385.5350 1120.0000 388.5350 ;
      RECT 1114.5000 383.4400 1120.0000 385.5350 ;
      RECT 1076.5000 383.4400 1111.5000 386.4400 ;
      RECT 1060.5000 383.4400 1073.5000 386.4400 ;
      RECT 1052.3500 383.4400 1057.5000 386.4400 ;
      RECT 1044.2000 383.4400 1049.3500 386.4400 ;
      RECT 1036.0500 383.4400 1041.2000 386.4400 ;
      RECT 1027.9000 383.4400 1033.0500 386.4400 ;
      RECT 1019.7500 383.4400 1024.9000 386.4400 ;
      RECT 1011.6000 383.4400 1016.7500 386.4400 ;
      RECT 1003.4500 383.4400 1008.6000 386.4400 ;
      RECT 995.3000 383.4400 1000.4500 386.4400 ;
      RECT 987.1500 383.4400 992.3000 386.4400 ;
      RECT 979.0000 383.4400 984.1500 386.4400 ;
      RECT 970.8500 383.4400 976.0000 386.4400 ;
      RECT 962.7000 383.4400 967.8500 386.4400 ;
      RECT 954.5500 383.4400 959.7000 386.4400 ;
      RECT 946.4000 383.4400 951.5500 386.4400 ;
      RECT 938.2500 383.4400 943.4000 386.4400 ;
      RECT 930.1000 383.4400 935.2500 386.4400 ;
      RECT 921.9500 383.4400 927.1000 386.4400 ;
      RECT 913.8000 383.4400 918.9500 386.4400 ;
      RECT 905.6500 383.4400 910.8000 386.4400 ;
      RECT 897.5000 383.4400 902.6500 386.4400 ;
      RECT 889.3500 383.4400 894.5000 386.4400 ;
      RECT 881.2000 383.4400 886.3500 386.4400 ;
      RECT 873.0500 383.4400 878.2000 386.4400 ;
      RECT 864.9000 383.4400 870.0500 386.4400 ;
      RECT 856.7500 383.4400 861.9000 386.4400 ;
      RECT 848.6000 383.4400 853.7500 386.4400 ;
      RECT 840.4500 383.4400 845.6000 386.4400 ;
      RECT 832.3000 383.4400 837.4500 386.4400 ;
      RECT 824.1500 383.4400 829.3000 386.4400 ;
      RECT 816.0000 383.4400 821.1500 386.4400 ;
      RECT 807.8500 383.4400 813.0000 386.4400 ;
      RECT 799.7000 383.4400 804.8500 386.4400 ;
      RECT 791.5500 383.4400 796.7000 386.4400 ;
      RECT 783.4000 383.4400 788.5500 386.4400 ;
      RECT 775.2500 383.4400 780.4000 386.4400 ;
      RECT 767.1000 383.4400 772.2500 386.4400 ;
      RECT 758.9500 383.4400 764.1000 386.4400 ;
      RECT 750.8000 383.4400 755.9500 386.4400 ;
      RECT 742.6500 383.4400 747.8000 386.4400 ;
      RECT 734.5000 383.4400 739.6500 386.4400 ;
      RECT 726.3500 383.4400 731.5000 386.4400 ;
      RECT 718.2000 383.4400 723.3500 386.4400 ;
      RECT 710.0500 383.4400 715.2000 386.4400 ;
      RECT 701.9000 383.4400 707.0500 386.4400 ;
      RECT 693.7500 383.4400 698.9000 386.4400 ;
      RECT 685.6000 383.4400 690.7500 386.4400 ;
      RECT 677.4500 383.4400 682.6000 386.4400 ;
      RECT 669.3000 383.4400 674.4500 386.4400 ;
      RECT 661.1500 383.4400 666.3000 386.4400 ;
      RECT 653.0000 383.4400 658.1500 386.4400 ;
      RECT 644.8500 383.4400 650.0000 386.4400 ;
      RECT 636.7000 383.4400 641.8500 386.4400 ;
      RECT 628.5500 383.4400 633.7000 386.4400 ;
      RECT 620.4000 383.4400 625.5500 386.4400 ;
      RECT 612.2500 383.4400 617.4000 386.4400 ;
      RECT 604.1000 383.4400 609.2500 386.4400 ;
      RECT 595.9500 383.4400 601.1000 386.4400 ;
      RECT 587.8000 383.4400 592.9500 386.4400 ;
      RECT 579.6500 383.4400 584.8000 386.4400 ;
      RECT 571.5000 383.4400 576.6500 386.4400 ;
      RECT 563.3500 383.4400 568.5000 386.4400 ;
      RECT 555.2000 383.4400 560.3500 386.4400 ;
      RECT 547.0500 383.4400 552.2000 386.4400 ;
      RECT 538.9000 383.4400 544.0500 386.4400 ;
      RECT 530.7500 383.4400 535.9000 386.4400 ;
      RECT 522.6000 383.4400 527.7500 386.4400 ;
      RECT 514.4500 383.4400 519.6000 386.4400 ;
      RECT 506.3000 383.4400 511.4500 386.4400 ;
      RECT 498.1500 383.4400 503.3000 386.4400 ;
      RECT 490.0000 383.4400 495.1500 386.4400 ;
      RECT 481.8500 383.4400 487.0000 386.4400 ;
      RECT 473.7000 383.4400 478.8500 386.4400 ;
      RECT 465.5500 383.4400 470.7000 386.4400 ;
      RECT 457.4000 383.4400 462.5500 386.4400 ;
      RECT 449.2500 383.4400 454.4000 386.4400 ;
      RECT 441.1000 383.4400 446.2500 386.4400 ;
      RECT 432.9500 383.4400 438.1000 386.4400 ;
      RECT 424.8000 383.4400 429.9500 386.4400 ;
      RECT 416.6500 383.4400 421.8000 386.4400 ;
      RECT 396.5000 383.4400 413.6500 386.4400 ;
      RECT 8.5000 383.4400 393.5000 386.4400 ;
      RECT 0.0000 383.4400 5.5000 386.4400 ;
      RECT 0.0000 381.4400 1120.0000 383.4400 ;
      RECT 0.0000 379.3450 1115.5000 381.4400 ;
      RECT 1118.5000 378.4400 1120.0000 381.4400 ;
      RECT 1114.5000 378.4400 1115.5000 379.3450 ;
      RECT 1114.5000 376.3450 1120.0000 378.4400 ;
      RECT 1076.5000 376.3450 1111.5000 379.3450 ;
      RECT 1060.5000 376.3450 1073.5000 379.3450 ;
      RECT 1052.3500 376.3450 1057.5000 379.3450 ;
      RECT 1044.2000 376.3450 1049.3500 379.3450 ;
      RECT 1036.0500 376.3450 1041.2000 379.3450 ;
      RECT 1027.9000 376.3450 1033.0500 379.3450 ;
      RECT 1019.7500 376.3450 1024.9000 379.3450 ;
      RECT 1011.6000 376.3450 1016.7500 379.3450 ;
      RECT 1003.4500 376.3450 1008.6000 379.3450 ;
      RECT 995.3000 376.3450 1000.4500 379.3450 ;
      RECT 987.1500 376.3450 992.3000 379.3450 ;
      RECT 979.0000 376.3450 984.1500 379.3450 ;
      RECT 970.8500 376.3450 976.0000 379.3450 ;
      RECT 962.7000 376.3450 967.8500 379.3450 ;
      RECT 954.5500 376.3450 959.7000 379.3450 ;
      RECT 946.4000 376.3450 951.5500 379.3450 ;
      RECT 938.2500 376.3450 943.4000 379.3450 ;
      RECT 930.1000 376.3450 935.2500 379.3450 ;
      RECT 921.9500 376.3450 927.1000 379.3450 ;
      RECT 913.8000 376.3450 918.9500 379.3450 ;
      RECT 905.6500 376.3450 910.8000 379.3450 ;
      RECT 897.5000 376.3450 902.6500 379.3450 ;
      RECT 889.3500 376.3450 894.5000 379.3450 ;
      RECT 881.2000 376.3450 886.3500 379.3450 ;
      RECT 873.0500 376.3450 878.2000 379.3450 ;
      RECT 864.9000 376.3450 870.0500 379.3450 ;
      RECT 856.7500 376.3450 861.9000 379.3450 ;
      RECT 848.6000 376.3450 853.7500 379.3450 ;
      RECT 840.4500 376.3450 845.6000 379.3450 ;
      RECT 832.3000 376.3450 837.4500 379.3450 ;
      RECT 824.1500 376.3450 829.3000 379.3450 ;
      RECT 816.0000 376.3450 821.1500 379.3450 ;
      RECT 807.8500 376.3450 813.0000 379.3450 ;
      RECT 799.7000 376.3450 804.8500 379.3450 ;
      RECT 791.5500 376.3450 796.7000 379.3450 ;
      RECT 783.4000 376.3450 788.5500 379.3450 ;
      RECT 775.2500 376.3450 780.4000 379.3450 ;
      RECT 767.1000 376.3450 772.2500 379.3450 ;
      RECT 758.9500 376.3450 764.1000 379.3450 ;
      RECT 750.8000 376.3450 755.9500 379.3450 ;
      RECT 742.6500 376.3450 747.8000 379.3450 ;
      RECT 734.5000 376.3450 739.6500 379.3450 ;
      RECT 726.3500 376.3450 731.5000 379.3450 ;
      RECT 718.2000 376.3450 723.3500 379.3450 ;
      RECT 710.0500 376.3450 715.2000 379.3450 ;
      RECT 701.9000 376.3450 707.0500 379.3450 ;
      RECT 693.7500 376.3450 698.9000 379.3450 ;
      RECT 685.6000 376.3450 690.7500 379.3450 ;
      RECT 677.4500 376.3450 682.6000 379.3450 ;
      RECT 669.3000 376.3450 674.4500 379.3450 ;
      RECT 661.1500 376.3450 666.3000 379.3450 ;
      RECT 653.0000 376.3450 658.1500 379.3450 ;
      RECT 644.8500 376.3450 650.0000 379.3450 ;
      RECT 636.7000 376.3450 641.8500 379.3450 ;
      RECT 628.5500 376.3450 633.7000 379.3450 ;
      RECT 620.4000 376.3450 625.5500 379.3450 ;
      RECT 612.2500 376.3450 617.4000 379.3450 ;
      RECT 604.1000 376.3450 609.2500 379.3450 ;
      RECT 595.9500 376.3450 601.1000 379.3450 ;
      RECT 587.8000 376.3450 592.9500 379.3450 ;
      RECT 579.6500 376.3450 584.8000 379.3450 ;
      RECT 571.5000 376.3450 576.6500 379.3450 ;
      RECT 563.3500 376.3450 568.5000 379.3450 ;
      RECT 555.2000 376.3450 560.3500 379.3450 ;
      RECT 547.0500 376.3450 552.2000 379.3450 ;
      RECT 538.9000 376.3450 544.0500 379.3450 ;
      RECT 530.7500 376.3450 535.9000 379.3450 ;
      RECT 522.6000 376.3450 527.7500 379.3450 ;
      RECT 514.4500 376.3450 519.6000 379.3450 ;
      RECT 506.3000 376.3450 511.4500 379.3450 ;
      RECT 498.1500 376.3450 503.3000 379.3450 ;
      RECT 490.0000 376.3450 495.1500 379.3450 ;
      RECT 481.8500 376.3450 487.0000 379.3450 ;
      RECT 473.7000 376.3450 478.8500 379.3450 ;
      RECT 465.5500 376.3450 470.7000 379.3450 ;
      RECT 457.4000 376.3450 462.5500 379.3450 ;
      RECT 449.2500 376.3450 454.4000 379.3450 ;
      RECT 441.1000 376.3450 446.2500 379.3450 ;
      RECT 432.9500 376.3450 438.1000 379.3450 ;
      RECT 424.8000 376.3450 429.9500 379.3450 ;
      RECT 416.6500 376.3450 421.8000 379.3450 ;
      RECT 396.5000 376.3450 413.6500 379.3450 ;
      RECT 8.5000 376.3450 393.5000 379.3450 ;
      RECT 0.0000 376.3450 5.5000 379.3450 ;
      RECT 0.0000 376.3000 1120.0000 376.3450 ;
      RECT 1073.5000 376.1000 1120.0000 376.3000 ;
      RECT 1116.6000 374.3450 1120.0000 376.1000 ;
      RECT 1073.5000 373.3000 1113.6000 376.1000 ;
      RECT 0.0000 373.3000 1070.5000 376.3000 ;
      RECT 0.0000 372.2500 1113.6000 373.3000 ;
      RECT 1118.5000 371.3450 1120.0000 374.3450 ;
      RECT 1114.5000 369.2500 1120.0000 371.3450 ;
      RECT 1076.5000 369.2500 1111.5000 372.2500 ;
      RECT 1060.5000 369.2500 1073.5000 372.2500 ;
      RECT 1052.3500 369.2500 1057.5000 372.2500 ;
      RECT 1044.2000 369.2500 1049.3500 372.2500 ;
      RECT 1036.0500 369.2500 1041.2000 372.2500 ;
      RECT 1027.9000 369.2500 1033.0500 372.2500 ;
      RECT 1019.7500 369.2500 1024.9000 372.2500 ;
      RECT 1011.6000 369.2500 1016.7500 372.2500 ;
      RECT 1003.4500 369.2500 1008.6000 372.2500 ;
      RECT 995.3000 369.2500 1000.4500 372.2500 ;
      RECT 987.1500 369.2500 992.3000 372.2500 ;
      RECT 979.0000 369.2500 984.1500 372.2500 ;
      RECT 970.8500 369.2500 976.0000 372.2500 ;
      RECT 962.7000 369.2500 967.8500 372.2500 ;
      RECT 954.5500 369.2500 959.7000 372.2500 ;
      RECT 946.4000 369.2500 951.5500 372.2500 ;
      RECT 938.2500 369.2500 943.4000 372.2500 ;
      RECT 930.1000 369.2500 935.2500 372.2500 ;
      RECT 921.9500 369.2500 927.1000 372.2500 ;
      RECT 913.8000 369.2500 918.9500 372.2500 ;
      RECT 905.6500 369.2500 910.8000 372.2500 ;
      RECT 897.5000 369.2500 902.6500 372.2500 ;
      RECT 889.3500 369.2500 894.5000 372.2500 ;
      RECT 881.2000 369.2500 886.3500 372.2500 ;
      RECT 873.0500 369.2500 878.2000 372.2500 ;
      RECT 864.9000 369.2500 870.0500 372.2500 ;
      RECT 856.7500 369.2500 861.9000 372.2500 ;
      RECT 848.6000 369.2500 853.7500 372.2500 ;
      RECT 840.4500 369.2500 845.6000 372.2500 ;
      RECT 832.3000 369.2500 837.4500 372.2500 ;
      RECT 824.1500 369.2500 829.3000 372.2500 ;
      RECT 816.0000 369.2500 821.1500 372.2500 ;
      RECT 807.8500 369.2500 813.0000 372.2500 ;
      RECT 799.7000 369.2500 804.8500 372.2500 ;
      RECT 791.5500 369.2500 796.7000 372.2500 ;
      RECT 783.4000 369.2500 788.5500 372.2500 ;
      RECT 775.2500 369.2500 780.4000 372.2500 ;
      RECT 767.1000 369.2500 772.2500 372.2500 ;
      RECT 758.9500 369.2500 764.1000 372.2500 ;
      RECT 750.8000 369.2500 755.9500 372.2500 ;
      RECT 742.6500 369.2500 747.8000 372.2500 ;
      RECT 734.5000 369.2500 739.6500 372.2500 ;
      RECT 726.3500 369.2500 731.5000 372.2500 ;
      RECT 718.2000 369.2500 723.3500 372.2500 ;
      RECT 710.0500 369.2500 715.2000 372.2500 ;
      RECT 701.9000 369.2500 707.0500 372.2500 ;
      RECT 693.7500 369.2500 698.9000 372.2500 ;
      RECT 685.6000 369.2500 690.7500 372.2500 ;
      RECT 677.4500 369.2500 682.6000 372.2500 ;
      RECT 669.3000 369.2500 674.4500 372.2500 ;
      RECT 661.1500 369.2500 666.3000 372.2500 ;
      RECT 653.0000 369.2500 658.1500 372.2500 ;
      RECT 644.8500 369.2500 650.0000 372.2500 ;
      RECT 636.7000 369.2500 641.8500 372.2500 ;
      RECT 628.5500 369.2500 633.7000 372.2500 ;
      RECT 620.4000 369.2500 625.5500 372.2500 ;
      RECT 612.2500 369.2500 617.4000 372.2500 ;
      RECT 604.1000 369.2500 609.2500 372.2500 ;
      RECT 595.9500 369.2500 601.1000 372.2500 ;
      RECT 587.8000 369.2500 592.9500 372.2500 ;
      RECT 579.6500 369.2500 584.8000 372.2500 ;
      RECT 571.5000 369.2500 576.6500 372.2500 ;
      RECT 563.3500 369.2500 568.5000 372.2500 ;
      RECT 555.2000 369.2500 560.3500 372.2500 ;
      RECT 547.0500 369.2500 552.2000 372.2500 ;
      RECT 538.9000 369.2500 544.0500 372.2500 ;
      RECT 530.7500 369.2500 535.9000 372.2500 ;
      RECT 522.6000 369.2500 527.7500 372.2500 ;
      RECT 514.4500 369.2500 519.6000 372.2500 ;
      RECT 506.3000 369.2500 511.4500 372.2500 ;
      RECT 498.1500 369.2500 503.3000 372.2500 ;
      RECT 490.0000 369.2500 495.1500 372.2500 ;
      RECT 481.8500 369.2500 487.0000 372.2500 ;
      RECT 473.7000 369.2500 478.8500 372.2500 ;
      RECT 465.5500 369.2500 470.7000 372.2500 ;
      RECT 457.4000 369.2500 462.5500 372.2500 ;
      RECT 449.2500 369.2500 454.4000 372.2500 ;
      RECT 441.1000 369.2500 446.2500 372.2500 ;
      RECT 432.9500 369.2500 438.1000 372.2500 ;
      RECT 424.8000 369.2500 429.9500 372.2500 ;
      RECT 416.6500 369.2500 421.8000 372.2500 ;
      RECT 396.5000 369.2500 413.6500 372.2500 ;
      RECT 8.5000 369.2500 393.5000 372.2500 ;
      RECT 0.0000 369.2500 5.5000 372.2500 ;
      RECT 0.0000 367.7000 1120.0000 369.2500 ;
      RECT 1116.6000 367.2500 1120.0000 367.7000 ;
      RECT 0.0000 365.1550 1113.6000 367.7000 ;
      RECT 1118.5000 364.2500 1120.0000 367.2500 ;
      RECT 1114.5000 362.1550 1120.0000 364.2500 ;
      RECT 1076.5000 362.1550 1111.5000 365.1550 ;
      RECT 1060.5000 362.1550 1073.5000 365.1550 ;
      RECT 1052.3500 362.1550 1057.5000 365.1550 ;
      RECT 1044.2000 362.1550 1049.3500 365.1550 ;
      RECT 1036.0500 362.1550 1041.2000 365.1550 ;
      RECT 1027.9000 362.1550 1033.0500 365.1550 ;
      RECT 1019.7500 362.1550 1024.9000 365.1550 ;
      RECT 1011.6000 362.1550 1016.7500 365.1550 ;
      RECT 1003.4500 362.1550 1008.6000 365.1550 ;
      RECT 995.3000 362.1550 1000.4500 365.1550 ;
      RECT 987.1500 362.1550 992.3000 365.1550 ;
      RECT 979.0000 362.1550 984.1500 365.1550 ;
      RECT 970.8500 362.1550 976.0000 365.1550 ;
      RECT 962.7000 362.1550 967.8500 365.1550 ;
      RECT 954.5500 362.1550 959.7000 365.1550 ;
      RECT 946.4000 362.1550 951.5500 365.1550 ;
      RECT 938.2500 362.1550 943.4000 365.1550 ;
      RECT 930.1000 362.1550 935.2500 365.1550 ;
      RECT 921.9500 362.1550 927.1000 365.1550 ;
      RECT 913.8000 362.1550 918.9500 365.1550 ;
      RECT 905.6500 362.1550 910.8000 365.1550 ;
      RECT 897.5000 362.1550 902.6500 365.1550 ;
      RECT 889.3500 362.1550 894.5000 365.1550 ;
      RECT 881.2000 362.1550 886.3500 365.1550 ;
      RECT 873.0500 362.1550 878.2000 365.1550 ;
      RECT 864.9000 362.1550 870.0500 365.1550 ;
      RECT 856.7500 362.1550 861.9000 365.1550 ;
      RECT 848.6000 362.1550 853.7500 365.1550 ;
      RECT 840.4500 362.1550 845.6000 365.1550 ;
      RECT 832.3000 362.1550 837.4500 365.1550 ;
      RECT 824.1500 362.1550 829.3000 365.1550 ;
      RECT 816.0000 362.1550 821.1500 365.1550 ;
      RECT 807.8500 362.1550 813.0000 365.1550 ;
      RECT 799.7000 362.1550 804.8500 365.1550 ;
      RECT 791.5500 362.1550 796.7000 365.1550 ;
      RECT 783.4000 362.1550 788.5500 365.1550 ;
      RECT 775.2500 362.1550 780.4000 365.1550 ;
      RECT 767.1000 362.1550 772.2500 365.1550 ;
      RECT 758.9500 362.1550 764.1000 365.1550 ;
      RECT 750.8000 362.1550 755.9500 365.1550 ;
      RECT 742.6500 362.1550 747.8000 365.1550 ;
      RECT 734.5000 362.1550 739.6500 365.1550 ;
      RECT 726.3500 362.1550 731.5000 365.1550 ;
      RECT 718.2000 362.1550 723.3500 365.1550 ;
      RECT 710.0500 362.1550 715.2000 365.1550 ;
      RECT 701.9000 362.1550 707.0500 365.1550 ;
      RECT 693.7500 362.1550 698.9000 365.1550 ;
      RECT 685.6000 362.1550 690.7500 365.1550 ;
      RECT 677.4500 362.1550 682.6000 365.1550 ;
      RECT 669.3000 362.1550 674.4500 365.1550 ;
      RECT 661.1500 362.1550 666.3000 365.1550 ;
      RECT 653.0000 362.1550 658.1500 365.1550 ;
      RECT 644.8500 362.1550 650.0000 365.1550 ;
      RECT 636.7000 362.1550 641.8500 365.1550 ;
      RECT 628.5500 362.1550 633.7000 365.1550 ;
      RECT 620.4000 362.1550 625.5500 365.1550 ;
      RECT 612.2500 362.1550 617.4000 365.1550 ;
      RECT 604.1000 362.1550 609.2500 365.1550 ;
      RECT 595.9500 362.1550 601.1000 365.1550 ;
      RECT 587.8000 362.1550 592.9500 365.1550 ;
      RECT 579.6500 362.1550 584.8000 365.1550 ;
      RECT 571.5000 362.1550 576.6500 365.1550 ;
      RECT 563.3500 362.1550 568.5000 365.1550 ;
      RECT 555.2000 362.1550 560.3500 365.1550 ;
      RECT 547.0500 362.1550 552.2000 365.1550 ;
      RECT 538.9000 362.1550 544.0500 365.1550 ;
      RECT 530.7500 362.1550 535.9000 365.1550 ;
      RECT 522.6000 362.1550 527.7500 365.1550 ;
      RECT 514.4500 362.1550 519.6000 365.1550 ;
      RECT 506.3000 362.1550 511.4500 365.1550 ;
      RECT 498.1500 362.1550 503.3000 365.1550 ;
      RECT 490.0000 362.1550 495.1500 365.1550 ;
      RECT 481.8500 362.1550 487.0000 365.1550 ;
      RECT 473.7000 362.1550 478.8500 365.1550 ;
      RECT 465.5500 362.1550 470.7000 365.1550 ;
      RECT 457.4000 362.1550 462.5500 365.1550 ;
      RECT 449.2500 362.1550 454.4000 365.1550 ;
      RECT 441.1000 362.1550 446.2500 365.1550 ;
      RECT 432.9500 362.1550 438.1000 365.1550 ;
      RECT 424.8000 362.1550 429.9500 365.1550 ;
      RECT 416.6500 362.1550 421.8000 365.1550 ;
      RECT 396.5000 362.1550 413.6500 365.1550 ;
      RECT 8.5000 362.1550 393.5000 365.1550 ;
      RECT 0.0000 362.1550 5.5000 365.1550 ;
      RECT 0.0000 360.7000 1120.0000 362.1550 ;
      RECT 1116.6000 360.1550 1120.0000 360.7000 ;
      RECT 0.0000 358.0600 1113.6000 360.7000 ;
      RECT 1118.5000 357.1550 1120.0000 360.1550 ;
      RECT 1114.5000 355.0600 1120.0000 357.1550 ;
      RECT 1076.5000 355.0600 1111.5000 358.0600 ;
      RECT 1060.5000 355.0600 1073.5000 358.0600 ;
      RECT 1052.3500 355.0600 1057.5000 358.0600 ;
      RECT 1044.2000 355.0600 1049.3500 358.0600 ;
      RECT 1036.0500 355.0600 1041.2000 358.0600 ;
      RECT 1027.9000 355.0600 1033.0500 358.0600 ;
      RECT 1019.7500 355.0600 1024.9000 358.0600 ;
      RECT 1011.6000 355.0600 1016.7500 358.0600 ;
      RECT 1003.4500 355.0600 1008.6000 358.0600 ;
      RECT 995.3000 355.0600 1000.4500 358.0600 ;
      RECT 987.1500 355.0600 992.3000 358.0600 ;
      RECT 979.0000 355.0600 984.1500 358.0600 ;
      RECT 970.8500 355.0600 976.0000 358.0600 ;
      RECT 962.7000 355.0600 967.8500 358.0600 ;
      RECT 954.5500 355.0600 959.7000 358.0600 ;
      RECT 946.4000 355.0600 951.5500 358.0600 ;
      RECT 938.2500 355.0600 943.4000 358.0600 ;
      RECT 930.1000 355.0600 935.2500 358.0600 ;
      RECT 921.9500 355.0600 927.1000 358.0600 ;
      RECT 913.8000 355.0600 918.9500 358.0600 ;
      RECT 905.6500 355.0600 910.8000 358.0600 ;
      RECT 897.5000 355.0600 902.6500 358.0600 ;
      RECT 889.3500 355.0600 894.5000 358.0600 ;
      RECT 881.2000 355.0600 886.3500 358.0600 ;
      RECT 873.0500 355.0600 878.2000 358.0600 ;
      RECT 864.9000 355.0600 870.0500 358.0600 ;
      RECT 856.7500 355.0600 861.9000 358.0600 ;
      RECT 848.6000 355.0600 853.7500 358.0600 ;
      RECT 840.4500 355.0600 845.6000 358.0600 ;
      RECT 832.3000 355.0600 837.4500 358.0600 ;
      RECT 824.1500 355.0600 829.3000 358.0600 ;
      RECT 816.0000 355.0600 821.1500 358.0600 ;
      RECT 807.8500 355.0600 813.0000 358.0600 ;
      RECT 799.7000 355.0600 804.8500 358.0600 ;
      RECT 791.5500 355.0600 796.7000 358.0600 ;
      RECT 783.4000 355.0600 788.5500 358.0600 ;
      RECT 775.2500 355.0600 780.4000 358.0600 ;
      RECT 767.1000 355.0600 772.2500 358.0600 ;
      RECT 758.9500 355.0600 764.1000 358.0600 ;
      RECT 750.8000 355.0600 755.9500 358.0600 ;
      RECT 742.6500 355.0600 747.8000 358.0600 ;
      RECT 734.5000 355.0600 739.6500 358.0600 ;
      RECT 726.3500 355.0600 731.5000 358.0600 ;
      RECT 718.2000 355.0600 723.3500 358.0600 ;
      RECT 710.0500 355.0600 715.2000 358.0600 ;
      RECT 701.9000 355.0600 707.0500 358.0600 ;
      RECT 693.7500 355.0600 698.9000 358.0600 ;
      RECT 685.6000 355.0600 690.7500 358.0600 ;
      RECT 677.4500 355.0600 682.6000 358.0600 ;
      RECT 669.3000 355.0600 674.4500 358.0600 ;
      RECT 661.1500 355.0600 666.3000 358.0600 ;
      RECT 653.0000 355.0600 658.1500 358.0600 ;
      RECT 644.8500 355.0600 650.0000 358.0600 ;
      RECT 636.7000 355.0600 641.8500 358.0600 ;
      RECT 628.5500 355.0600 633.7000 358.0600 ;
      RECT 620.4000 355.0600 625.5500 358.0600 ;
      RECT 612.2500 355.0600 617.4000 358.0600 ;
      RECT 604.1000 355.0600 609.2500 358.0600 ;
      RECT 595.9500 355.0600 601.1000 358.0600 ;
      RECT 587.8000 355.0600 592.9500 358.0600 ;
      RECT 579.6500 355.0600 584.8000 358.0600 ;
      RECT 571.5000 355.0600 576.6500 358.0600 ;
      RECT 563.3500 355.0600 568.5000 358.0600 ;
      RECT 555.2000 355.0600 560.3500 358.0600 ;
      RECT 547.0500 355.0600 552.2000 358.0600 ;
      RECT 538.9000 355.0600 544.0500 358.0600 ;
      RECT 530.7500 355.0600 535.9000 358.0600 ;
      RECT 522.6000 355.0600 527.7500 358.0600 ;
      RECT 514.4500 355.0600 519.6000 358.0600 ;
      RECT 506.3000 355.0600 511.4500 358.0600 ;
      RECT 498.1500 355.0600 503.3000 358.0600 ;
      RECT 490.0000 355.0600 495.1500 358.0600 ;
      RECT 481.8500 355.0600 487.0000 358.0600 ;
      RECT 473.7000 355.0600 478.8500 358.0600 ;
      RECT 465.5500 355.0600 470.7000 358.0600 ;
      RECT 457.4000 355.0600 462.5500 358.0600 ;
      RECT 449.2500 355.0600 454.4000 358.0600 ;
      RECT 441.1000 355.0600 446.2500 358.0600 ;
      RECT 432.9500 355.0600 438.1000 358.0600 ;
      RECT 424.8000 355.0600 429.9500 358.0600 ;
      RECT 416.6500 355.0600 421.8000 358.0600 ;
      RECT 396.5000 355.0600 413.6500 358.0600 ;
      RECT 8.5000 355.0600 393.5000 358.0600 ;
      RECT 0.0000 355.0600 5.5000 358.0600 ;
      RECT 0.0000 353.5000 1120.0000 355.0600 ;
      RECT 1116.6000 353.0600 1120.0000 353.5000 ;
      RECT 0.0000 350.9650 1113.6000 353.5000 ;
      RECT 1118.5000 350.0600 1120.0000 353.0600 ;
      RECT 1114.5000 347.9650 1120.0000 350.0600 ;
      RECT 1076.5000 347.9650 1111.5000 350.9650 ;
      RECT 1060.5000 347.9650 1073.5000 350.9650 ;
      RECT 1052.3500 347.9650 1057.5000 350.9650 ;
      RECT 1044.2000 347.9650 1049.3500 350.9650 ;
      RECT 1036.0500 347.9650 1041.2000 350.9650 ;
      RECT 1027.9000 347.9650 1033.0500 350.9650 ;
      RECT 1019.7500 347.9650 1024.9000 350.9650 ;
      RECT 1011.6000 347.9650 1016.7500 350.9650 ;
      RECT 1003.4500 347.9650 1008.6000 350.9650 ;
      RECT 995.3000 347.9650 1000.4500 350.9650 ;
      RECT 987.1500 347.9650 992.3000 350.9650 ;
      RECT 979.0000 347.9650 984.1500 350.9650 ;
      RECT 970.8500 347.9650 976.0000 350.9650 ;
      RECT 962.7000 347.9650 967.8500 350.9650 ;
      RECT 954.5500 347.9650 959.7000 350.9650 ;
      RECT 946.4000 347.9650 951.5500 350.9650 ;
      RECT 938.2500 347.9650 943.4000 350.9650 ;
      RECT 930.1000 347.9650 935.2500 350.9650 ;
      RECT 921.9500 347.9650 927.1000 350.9650 ;
      RECT 913.8000 347.9650 918.9500 350.9650 ;
      RECT 905.6500 347.9650 910.8000 350.9650 ;
      RECT 897.5000 347.9650 902.6500 350.9650 ;
      RECT 889.3500 347.9650 894.5000 350.9650 ;
      RECT 881.2000 347.9650 886.3500 350.9650 ;
      RECT 873.0500 347.9650 878.2000 350.9650 ;
      RECT 864.9000 347.9650 870.0500 350.9650 ;
      RECT 856.7500 347.9650 861.9000 350.9650 ;
      RECT 848.6000 347.9650 853.7500 350.9650 ;
      RECT 840.4500 347.9650 845.6000 350.9650 ;
      RECT 832.3000 347.9650 837.4500 350.9650 ;
      RECT 824.1500 347.9650 829.3000 350.9650 ;
      RECT 816.0000 347.9650 821.1500 350.9650 ;
      RECT 807.8500 347.9650 813.0000 350.9650 ;
      RECT 799.7000 347.9650 804.8500 350.9650 ;
      RECT 791.5500 347.9650 796.7000 350.9650 ;
      RECT 783.4000 347.9650 788.5500 350.9650 ;
      RECT 775.2500 347.9650 780.4000 350.9650 ;
      RECT 767.1000 347.9650 772.2500 350.9650 ;
      RECT 758.9500 347.9650 764.1000 350.9650 ;
      RECT 750.8000 347.9650 755.9500 350.9650 ;
      RECT 742.6500 347.9650 747.8000 350.9650 ;
      RECT 734.5000 347.9650 739.6500 350.9650 ;
      RECT 726.3500 347.9650 731.5000 350.9650 ;
      RECT 718.2000 347.9650 723.3500 350.9650 ;
      RECT 710.0500 347.9650 715.2000 350.9650 ;
      RECT 701.9000 347.9650 707.0500 350.9650 ;
      RECT 693.7500 347.9650 698.9000 350.9650 ;
      RECT 685.6000 347.9650 690.7500 350.9650 ;
      RECT 677.4500 347.9650 682.6000 350.9650 ;
      RECT 669.3000 347.9650 674.4500 350.9650 ;
      RECT 661.1500 347.9650 666.3000 350.9650 ;
      RECT 653.0000 347.9650 658.1500 350.9650 ;
      RECT 644.8500 347.9650 650.0000 350.9650 ;
      RECT 636.7000 347.9650 641.8500 350.9650 ;
      RECT 628.5500 347.9650 633.7000 350.9650 ;
      RECT 620.4000 347.9650 625.5500 350.9650 ;
      RECT 612.2500 347.9650 617.4000 350.9650 ;
      RECT 604.1000 347.9650 609.2500 350.9650 ;
      RECT 595.9500 347.9650 601.1000 350.9650 ;
      RECT 587.8000 347.9650 592.9500 350.9650 ;
      RECT 579.6500 347.9650 584.8000 350.9650 ;
      RECT 571.5000 347.9650 576.6500 350.9650 ;
      RECT 563.3500 347.9650 568.5000 350.9650 ;
      RECT 555.2000 347.9650 560.3500 350.9650 ;
      RECT 547.0500 347.9650 552.2000 350.9650 ;
      RECT 538.9000 347.9650 544.0500 350.9650 ;
      RECT 530.7500 347.9650 535.9000 350.9650 ;
      RECT 522.6000 347.9650 527.7500 350.9650 ;
      RECT 514.4500 347.9650 519.6000 350.9650 ;
      RECT 506.3000 347.9650 511.4500 350.9650 ;
      RECT 498.1500 347.9650 503.3000 350.9650 ;
      RECT 490.0000 347.9650 495.1500 350.9650 ;
      RECT 481.8500 347.9650 487.0000 350.9650 ;
      RECT 473.7000 347.9650 478.8500 350.9650 ;
      RECT 465.5500 347.9650 470.7000 350.9650 ;
      RECT 457.4000 347.9650 462.5500 350.9650 ;
      RECT 449.2500 347.9650 454.4000 350.9650 ;
      RECT 441.1000 347.9650 446.2500 350.9650 ;
      RECT 432.9500 347.9650 438.1000 350.9650 ;
      RECT 424.8000 347.9650 429.9500 350.9650 ;
      RECT 416.6500 347.9650 421.8000 350.9650 ;
      RECT 396.5000 347.9650 413.6500 350.9650 ;
      RECT 8.5000 347.9650 393.5000 350.9650 ;
      RECT 0.0000 347.9650 5.5000 350.9650 ;
      RECT 0.0000 346.5000 1120.0000 347.9650 ;
      RECT 1116.6000 345.9650 1120.0000 346.5000 ;
      RECT 0.0000 343.8700 1113.6000 346.5000 ;
      RECT 1118.5000 342.9650 1120.0000 345.9650 ;
      RECT 1114.5000 340.8700 1120.0000 342.9650 ;
      RECT 1076.5000 340.8700 1111.5000 343.8700 ;
      RECT 1060.5000 340.8700 1073.5000 343.8700 ;
      RECT 1052.3500 340.8700 1057.5000 343.8700 ;
      RECT 1044.2000 340.8700 1049.3500 343.8700 ;
      RECT 1036.0500 340.8700 1041.2000 343.8700 ;
      RECT 1027.9000 340.8700 1033.0500 343.8700 ;
      RECT 1019.7500 340.8700 1024.9000 343.8700 ;
      RECT 1011.6000 340.8700 1016.7500 343.8700 ;
      RECT 1003.4500 340.8700 1008.6000 343.8700 ;
      RECT 995.3000 340.8700 1000.4500 343.8700 ;
      RECT 987.1500 340.8700 992.3000 343.8700 ;
      RECT 979.0000 340.8700 984.1500 343.8700 ;
      RECT 970.8500 340.8700 976.0000 343.8700 ;
      RECT 962.7000 340.8700 967.8500 343.8700 ;
      RECT 954.5500 340.8700 959.7000 343.8700 ;
      RECT 946.4000 340.8700 951.5500 343.8700 ;
      RECT 938.2500 340.8700 943.4000 343.8700 ;
      RECT 930.1000 340.8700 935.2500 343.8700 ;
      RECT 921.9500 340.8700 927.1000 343.8700 ;
      RECT 913.8000 340.8700 918.9500 343.8700 ;
      RECT 905.6500 340.8700 910.8000 343.8700 ;
      RECT 897.5000 340.8700 902.6500 343.8700 ;
      RECT 889.3500 340.8700 894.5000 343.8700 ;
      RECT 881.2000 340.8700 886.3500 343.8700 ;
      RECT 873.0500 340.8700 878.2000 343.8700 ;
      RECT 864.9000 340.8700 870.0500 343.8700 ;
      RECT 856.7500 340.8700 861.9000 343.8700 ;
      RECT 848.6000 340.8700 853.7500 343.8700 ;
      RECT 840.4500 340.8700 845.6000 343.8700 ;
      RECT 832.3000 340.8700 837.4500 343.8700 ;
      RECT 824.1500 340.8700 829.3000 343.8700 ;
      RECT 816.0000 340.8700 821.1500 343.8700 ;
      RECT 807.8500 340.8700 813.0000 343.8700 ;
      RECT 799.7000 340.8700 804.8500 343.8700 ;
      RECT 791.5500 340.8700 796.7000 343.8700 ;
      RECT 783.4000 340.8700 788.5500 343.8700 ;
      RECT 775.2500 340.8700 780.4000 343.8700 ;
      RECT 767.1000 340.8700 772.2500 343.8700 ;
      RECT 758.9500 340.8700 764.1000 343.8700 ;
      RECT 750.8000 340.8700 755.9500 343.8700 ;
      RECT 742.6500 340.8700 747.8000 343.8700 ;
      RECT 734.5000 340.8700 739.6500 343.8700 ;
      RECT 726.3500 340.8700 731.5000 343.8700 ;
      RECT 718.2000 340.8700 723.3500 343.8700 ;
      RECT 710.0500 340.8700 715.2000 343.8700 ;
      RECT 701.9000 340.8700 707.0500 343.8700 ;
      RECT 693.7500 340.8700 698.9000 343.8700 ;
      RECT 685.6000 340.8700 690.7500 343.8700 ;
      RECT 677.4500 340.8700 682.6000 343.8700 ;
      RECT 669.3000 340.8700 674.4500 343.8700 ;
      RECT 661.1500 340.8700 666.3000 343.8700 ;
      RECT 653.0000 340.8700 658.1500 343.8700 ;
      RECT 644.8500 340.8700 650.0000 343.8700 ;
      RECT 636.7000 340.8700 641.8500 343.8700 ;
      RECT 628.5500 340.8700 633.7000 343.8700 ;
      RECT 620.4000 340.8700 625.5500 343.8700 ;
      RECT 612.2500 340.8700 617.4000 343.8700 ;
      RECT 604.1000 340.8700 609.2500 343.8700 ;
      RECT 595.9500 340.8700 601.1000 343.8700 ;
      RECT 587.8000 340.8700 592.9500 343.8700 ;
      RECT 579.6500 340.8700 584.8000 343.8700 ;
      RECT 571.5000 340.8700 576.6500 343.8700 ;
      RECT 563.3500 340.8700 568.5000 343.8700 ;
      RECT 555.2000 340.8700 560.3500 343.8700 ;
      RECT 547.0500 340.8700 552.2000 343.8700 ;
      RECT 538.9000 340.8700 544.0500 343.8700 ;
      RECT 530.7500 340.8700 535.9000 343.8700 ;
      RECT 522.6000 340.8700 527.7500 343.8700 ;
      RECT 514.4500 340.8700 519.6000 343.8700 ;
      RECT 506.3000 340.8700 511.4500 343.8700 ;
      RECT 498.1500 340.8700 503.3000 343.8700 ;
      RECT 490.0000 340.8700 495.1500 343.8700 ;
      RECT 481.8500 340.8700 487.0000 343.8700 ;
      RECT 473.7000 340.8700 478.8500 343.8700 ;
      RECT 465.5500 340.8700 470.7000 343.8700 ;
      RECT 457.4000 340.8700 462.5500 343.8700 ;
      RECT 449.2500 340.8700 454.4000 343.8700 ;
      RECT 441.1000 340.8700 446.2500 343.8700 ;
      RECT 432.9500 340.8700 438.1000 343.8700 ;
      RECT 424.8000 340.8700 429.9500 343.8700 ;
      RECT 416.6500 340.8700 421.8000 343.8700 ;
      RECT 396.5000 340.8700 413.6500 343.8700 ;
      RECT 346.5000 340.8700 393.5000 343.8700 ;
      RECT 46.5000 340.8700 343.5000 343.8700 ;
      RECT 8.5000 340.8700 43.5000 343.8700 ;
      RECT 0.0000 340.8700 5.5000 343.8700 ;
      RECT 0.0000 339.3000 1120.0000 340.8700 ;
      RECT 1116.6000 338.8700 1120.0000 339.3000 ;
      RECT 0.0000 336.7750 1113.6000 339.3000 ;
      RECT 1118.5000 335.8700 1120.0000 338.8700 ;
      RECT 1114.5000 333.7750 1120.0000 335.8700 ;
      RECT 1076.5000 333.7750 1111.5000 336.7750 ;
      RECT 1060.5000 333.7750 1073.5000 336.7750 ;
      RECT 1052.3500 333.7750 1057.5000 336.7750 ;
      RECT 1044.2000 333.7750 1049.3500 336.7750 ;
      RECT 1036.0500 333.7750 1041.2000 336.7750 ;
      RECT 1027.9000 333.7750 1033.0500 336.7750 ;
      RECT 1019.7500 333.7750 1024.9000 336.7750 ;
      RECT 1011.6000 333.7750 1016.7500 336.7750 ;
      RECT 1003.4500 333.7750 1008.6000 336.7750 ;
      RECT 995.3000 333.7750 1000.4500 336.7750 ;
      RECT 987.1500 333.7750 992.3000 336.7750 ;
      RECT 979.0000 333.7750 984.1500 336.7750 ;
      RECT 970.8500 333.7750 976.0000 336.7750 ;
      RECT 962.7000 333.7750 967.8500 336.7750 ;
      RECT 954.5500 333.7750 959.7000 336.7750 ;
      RECT 946.4000 333.7750 951.5500 336.7750 ;
      RECT 938.2500 333.7750 943.4000 336.7750 ;
      RECT 930.1000 333.7750 935.2500 336.7750 ;
      RECT 921.9500 333.7750 927.1000 336.7750 ;
      RECT 913.8000 333.7750 918.9500 336.7750 ;
      RECT 905.6500 333.7750 910.8000 336.7750 ;
      RECT 897.5000 333.7750 902.6500 336.7750 ;
      RECT 889.3500 333.7750 894.5000 336.7750 ;
      RECT 881.2000 333.7750 886.3500 336.7750 ;
      RECT 873.0500 333.7750 878.2000 336.7750 ;
      RECT 864.9000 333.7750 870.0500 336.7750 ;
      RECT 856.7500 333.7750 861.9000 336.7750 ;
      RECT 848.6000 333.7750 853.7500 336.7750 ;
      RECT 840.4500 333.7750 845.6000 336.7750 ;
      RECT 832.3000 333.7750 837.4500 336.7750 ;
      RECT 824.1500 333.7750 829.3000 336.7750 ;
      RECT 816.0000 333.7750 821.1500 336.7750 ;
      RECT 807.8500 333.7750 813.0000 336.7750 ;
      RECT 799.7000 333.7750 804.8500 336.7750 ;
      RECT 791.5500 333.7750 796.7000 336.7750 ;
      RECT 783.4000 333.7750 788.5500 336.7750 ;
      RECT 775.2500 333.7750 780.4000 336.7750 ;
      RECT 767.1000 333.7750 772.2500 336.7750 ;
      RECT 758.9500 333.7750 764.1000 336.7750 ;
      RECT 750.8000 333.7750 755.9500 336.7750 ;
      RECT 742.6500 333.7750 747.8000 336.7750 ;
      RECT 734.5000 333.7750 739.6500 336.7750 ;
      RECT 726.3500 333.7750 731.5000 336.7750 ;
      RECT 718.2000 333.7750 723.3500 336.7750 ;
      RECT 710.0500 333.7750 715.2000 336.7750 ;
      RECT 701.9000 333.7750 707.0500 336.7750 ;
      RECT 693.7500 333.7750 698.9000 336.7750 ;
      RECT 685.6000 333.7750 690.7500 336.7750 ;
      RECT 677.4500 333.7750 682.6000 336.7750 ;
      RECT 669.3000 333.7750 674.4500 336.7750 ;
      RECT 661.1500 333.7750 666.3000 336.7750 ;
      RECT 653.0000 333.7750 658.1500 336.7750 ;
      RECT 644.8500 333.7750 650.0000 336.7750 ;
      RECT 636.7000 333.7750 641.8500 336.7750 ;
      RECT 628.5500 333.7750 633.7000 336.7750 ;
      RECT 620.4000 333.7750 625.5500 336.7750 ;
      RECT 612.2500 333.7750 617.4000 336.7750 ;
      RECT 604.1000 333.7750 609.2500 336.7750 ;
      RECT 595.9500 333.7750 601.1000 336.7750 ;
      RECT 587.8000 333.7750 592.9500 336.7750 ;
      RECT 579.6500 333.7750 584.8000 336.7750 ;
      RECT 571.5000 333.7750 576.6500 336.7750 ;
      RECT 563.3500 333.7750 568.5000 336.7750 ;
      RECT 555.2000 333.7750 560.3500 336.7750 ;
      RECT 547.0500 333.7750 552.2000 336.7750 ;
      RECT 538.9000 333.7750 544.0500 336.7750 ;
      RECT 530.7500 333.7750 535.9000 336.7750 ;
      RECT 522.6000 333.7750 527.7500 336.7750 ;
      RECT 514.4500 333.7750 519.6000 336.7750 ;
      RECT 506.3000 333.7750 511.4500 336.7750 ;
      RECT 498.1500 333.7750 503.3000 336.7750 ;
      RECT 490.0000 333.7750 495.1500 336.7750 ;
      RECT 481.8500 333.7750 487.0000 336.7750 ;
      RECT 473.7000 333.7750 478.8500 336.7750 ;
      RECT 465.5500 333.7750 470.7000 336.7750 ;
      RECT 457.4000 333.7750 462.5500 336.7750 ;
      RECT 449.2500 333.7750 454.4000 336.7750 ;
      RECT 441.1000 333.7750 446.2500 336.7750 ;
      RECT 432.9500 333.7750 438.1000 336.7750 ;
      RECT 424.8000 333.7750 429.9500 336.7750 ;
      RECT 416.6500 333.7750 421.8000 336.7750 ;
      RECT 396.5000 333.7750 413.6500 336.7750 ;
      RECT 346.5000 333.7750 393.5000 336.7750 ;
      RECT 46.5000 333.7750 343.5000 336.7750 ;
      RECT 8.5000 333.7750 43.5000 336.7750 ;
      RECT 0.0000 333.7750 5.5000 336.7750 ;
      RECT 0.0000 332.3000 1120.0000 333.7750 ;
      RECT 1116.6000 331.7750 1120.0000 332.3000 ;
      RECT 0.0000 329.6800 1113.6000 332.3000 ;
      RECT 1118.5000 328.7750 1120.0000 331.7750 ;
      RECT 1114.5000 326.6800 1120.0000 328.7750 ;
      RECT 1076.5000 326.6800 1111.5000 329.6800 ;
      RECT 1060.5000 326.6800 1073.5000 329.6800 ;
      RECT 1052.3500 326.6800 1057.5000 329.6800 ;
      RECT 1044.2000 326.6800 1049.3500 329.6800 ;
      RECT 1036.0500 326.6800 1041.2000 329.6800 ;
      RECT 1027.9000 326.6800 1033.0500 329.6800 ;
      RECT 1019.7500 326.6800 1024.9000 329.6800 ;
      RECT 1011.6000 326.6800 1016.7500 329.6800 ;
      RECT 1003.4500 326.6800 1008.6000 329.6800 ;
      RECT 995.3000 326.6800 1000.4500 329.6800 ;
      RECT 987.1500 326.6800 992.3000 329.6800 ;
      RECT 979.0000 326.6800 984.1500 329.6800 ;
      RECT 970.8500 326.6800 976.0000 329.6800 ;
      RECT 962.7000 326.6800 967.8500 329.6800 ;
      RECT 954.5500 326.6800 959.7000 329.6800 ;
      RECT 946.4000 326.6800 951.5500 329.6800 ;
      RECT 938.2500 326.6800 943.4000 329.6800 ;
      RECT 930.1000 326.6800 935.2500 329.6800 ;
      RECT 921.9500 326.6800 927.1000 329.6800 ;
      RECT 913.8000 326.6800 918.9500 329.6800 ;
      RECT 905.6500 326.6800 910.8000 329.6800 ;
      RECT 897.5000 326.6800 902.6500 329.6800 ;
      RECT 889.3500 326.6800 894.5000 329.6800 ;
      RECT 881.2000 326.6800 886.3500 329.6800 ;
      RECT 873.0500 326.6800 878.2000 329.6800 ;
      RECT 864.9000 326.6800 870.0500 329.6800 ;
      RECT 856.7500 326.6800 861.9000 329.6800 ;
      RECT 848.6000 326.6800 853.7500 329.6800 ;
      RECT 840.4500 326.6800 845.6000 329.6800 ;
      RECT 832.3000 326.6800 837.4500 329.6800 ;
      RECT 824.1500 326.6800 829.3000 329.6800 ;
      RECT 816.0000 326.6800 821.1500 329.6800 ;
      RECT 807.8500 326.6800 813.0000 329.6800 ;
      RECT 799.7000 326.6800 804.8500 329.6800 ;
      RECT 791.5500 326.6800 796.7000 329.6800 ;
      RECT 783.4000 326.6800 788.5500 329.6800 ;
      RECT 775.2500 326.6800 780.4000 329.6800 ;
      RECT 767.1000 326.6800 772.2500 329.6800 ;
      RECT 758.9500 326.6800 764.1000 329.6800 ;
      RECT 750.8000 326.6800 755.9500 329.6800 ;
      RECT 742.6500 326.6800 747.8000 329.6800 ;
      RECT 734.5000 326.6800 739.6500 329.6800 ;
      RECT 726.3500 326.6800 731.5000 329.6800 ;
      RECT 718.2000 326.6800 723.3500 329.6800 ;
      RECT 710.0500 326.6800 715.2000 329.6800 ;
      RECT 701.9000 326.6800 707.0500 329.6800 ;
      RECT 693.7500 326.6800 698.9000 329.6800 ;
      RECT 685.6000 326.6800 690.7500 329.6800 ;
      RECT 677.4500 326.6800 682.6000 329.6800 ;
      RECT 669.3000 326.6800 674.4500 329.6800 ;
      RECT 661.1500 326.6800 666.3000 329.6800 ;
      RECT 653.0000 326.6800 658.1500 329.6800 ;
      RECT 644.8500 326.6800 650.0000 329.6800 ;
      RECT 636.7000 326.6800 641.8500 329.6800 ;
      RECT 628.5500 326.6800 633.7000 329.6800 ;
      RECT 620.4000 326.6800 625.5500 329.6800 ;
      RECT 612.2500 326.6800 617.4000 329.6800 ;
      RECT 604.1000 326.6800 609.2500 329.6800 ;
      RECT 595.9500 326.6800 601.1000 329.6800 ;
      RECT 587.8000 326.6800 592.9500 329.6800 ;
      RECT 579.6500 326.6800 584.8000 329.6800 ;
      RECT 571.5000 326.6800 576.6500 329.6800 ;
      RECT 563.3500 326.6800 568.5000 329.6800 ;
      RECT 555.2000 326.6800 560.3500 329.6800 ;
      RECT 547.0500 326.6800 552.2000 329.6800 ;
      RECT 538.9000 326.6800 544.0500 329.6800 ;
      RECT 530.7500 326.6800 535.9000 329.6800 ;
      RECT 522.6000 326.6800 527.7500 329.6800 ;
      RECT 514.4500 326.6800 519.6000 329.6800 ;
      RECT 506.3000 326.6800 511.4500 329.6800 ;
      RECT 498.1500 326.6800 503.3000 329.6800 ;
      RECT 490.0000 326.6800 495.1500 329.6800 ;
      RECT 481.8500 326.6800 487.0000 329.6800 ;
      RECT 473.7000 326.6800 478.8500 329.6800 ;
      RECT 465.5500 326.6800 470.7000 329.6800 ;
      RECT 457.4000 326.6800 462.5500 329.6800 ;
      RECT 449.2500 326.6800 454.4000 329.6800 ;
      RECT 441.1000 326.6800 446.2500 329.6800 ;
      RECT 432.9500 326.6800 438.1000 329.6800 ;
      RECT 424.8000 326.6800 429.9500 329.6800 ;
      RECT 416.6500 326.6800 421.8000 329.6800 ;
      RECT 396.5000 326.6800 413.6500 329.6800 ;
      RECT 346.5000 326.6800 393.5000 329.6800 ;
      RECT 326.4650 326.6800 343.5000 329.6800 ;
      RECT 317.9500 326.6800 323.4650 329.6800 ;
      RECT 309.4350 326.6800 314.9500 329.6800 ;
      RECT 300.9200 326.6800 306.4350 329.6800 ;
      RECT 292.4050 326.6800 297.9200 329.6800 ;
      RECT 283.8900 326.6800 289.4050 329.6800 ;
      RECT 275.3750 326.6800 280.8900 329.6800 ;
      RECT 266.8600 326.6800 272.3750 329.6800 ;
      RECT 258.3450 326.6800 263.8600 329.6800 ;
      RECT 249.8300 326.6800 255.3450 329.6800 ;
      RECT 241.3150 326.6800 246.8300 329.6800 ;
      RECT 232.8000 326.6800 238.3150 329.6800 ;
      RECT 224.2850 326.6800 229.8000 329.6800 ;
      RECT 215.7700 326.6800 221.2850 329.6800 ;
      RECT 207.2550 326.6800 212.7700 329.6800 ;
      RECT 198.7400 326.6800 204.2550 329.6800 ;
      RECT 190.2250 326.6800 195.7400 329.6800 ;
      RECT 181.7100 326.6800 187.2250 329.6800 ;
      RECT 173.1950 326.6800 178.7100 329.6800 ;
      RECT 164.6800 326.6800 170.1950 329.6800 ;
      RECT 156.1650 326.6800 161.6800 329.6800 ;
      RECT 147.6500 326.6800 153.1650 329.6800 ;
      RECT 139.1350 326.6800 144.6500 329.6800 ;
      RECT 130.6200 326.6800 136.1350 329.6800 ;
      RECT 122.1050 326.6800 127.6200 329.6800 ;
      RECT 113.5900 326.6800 119.1050 329.6800 ;
      RECT 105.0750 326.6800 110.5900 329.6800 ;
      RECT 96.5600 326.6800 102.0750 329.6800 ;
      RECT 88.0450 326.6800 93.5600 329.6800 ;
      RECT 79.5300 326.6800 85.0450 329.6800 ;
      RECT 71.0150 326.6800 76.5300 329.6800 ;
      RECT 62.5000 326.6800 68.0150 329.6800 ;
      RECT 46.5000 326.6800 59.5000 329.6800 ;
      RECT 8.5000 326.6800 43.5000 329.6800 ;
      RECT 0.0000 326.6800 5.5000 329.6800 ;
      RECT 0.0000 325.1000 1120.0000 326.6800 ;
      RECT 1116.6000 324.6800 1120.0000 325.1000 ;
      RECT 0.0000 322.5850 1113.6000 325.1000 ;
      RECT 1118.5000 321.6800 1120.0000 324.6800 ;
      RECT 1114.5000 319.5850 1120.0000 321.6800 ;
      RECT 1076.5000 319.5850 1111.5000 322.5850 ;
      RECT 1060.5000 319.5850 1073.5000 322.5850 ;
      RECT 1052.3500 319.5850 1057.5000 322.5850 ;
      RECT 1044.2000 319.5850 1049.3500 322.5850 ;
      RECT 1036.0500 319.5850 1041.2000 322.5850 ;
      RECT 1027.9000 319.5850 1033.0500 322.5850 ;
      RECT 1019.7500 319.5850 1024.9000 322.5850 ;
      RECT 1011.6000 319.5850 1016.7500 322.5850 ;
      RECT 1003.4500 319.5850 1008.6000 322.5850 ;
      RECT 995.3000 319.5850 1000.4500 322.5850 ;
      RECT 987.1500 319.5850 992.3000 322.5850 ;
      RECT 979.0000 319.5850 984.1500 322.5850 ;
      RECT 970.8500 319.5850 976.0000 322.5850 ;
      RECT 962.7000 319.5850 967.8500 322.5850 ;
      RECT 954.5500 319.5850 959.7000 322.5850 ;
      RECT 946.4000 319.5850 951.5500 322.5850 ;
      RECT 938.2500 319.5850 943.4000 322.5850 ;
      RECT 930.1000 319.5850 935.2500 322.5850 ;
      RECT 921.9500 319.5850 927.1000 322.5850 ;
      RECT 913.8000 319.5850 918.9500 322.5850 ;
      RECT 905.6500 319.5850 910.8000 322.5850 ;
      RECT 897.5000 319.5850 902.6500 322.5850 ;
      RECT 889.3500 319.5850 894.5000 322.5850 ;
      RECT 881.2000 319.5850 886.3500 322.5850 ;
      RECT 873.0500 319.5850 878.2000 322.5850 ;
      RECT 864.9000 319.5850 870.0500 322.5850 ;
      RECT 856.7500 319.5850 861.9000 322.5850 ;
      RECT 848.6000 319.5850 853.7500 322.5850 ;
      RECT 840.4500 319.5850 845.6000 322.5850 ;
      RECT 832.3000 319.5850 837.4500 322.5850 ;
      RECT 824.1500 319.5850 829.3000 322.5850 ;
      RECT 816.0000 319.5850 821.1500 322.5850 ;
      RECT 807.8500 319.5850 813.0000 322.5850 ;
      RECT 799.7000 319.5850 804.8500 322.5850 ;
      RECT 791.5500 319.5850 796.7000 322.5850 ;
      RECT 783.4000 319.5850 788.5500 322.5850 ;
      RECT 775.2500 319.5850 780.4000 322.5850 ;
      RECT 767.1000 319.5850 772.2500 322.5850 ;
      RECT 758.9500 319.5850 764.1000 322.5850 ;
      RECT 750.8000 319.5850 755.9500 322.5850 ;
      RECT 742.6500 319.5850 747.8000 322.5850 ;
      RECT 734.5000 319.5850 739.6500 322.5850 ;
      RECT 726.3500 319.5850 731.5000 322.5850 ;
      RECT 718.2000 319.5850 723.3500 322.5850 ;
      RECT 710.0500 319.5850 715.2000 322.5850 ;
      RECT 701.9000 319.5850 707.0500 322.5850 ;
      RECT 693.7500 319.5850 698.9000 322.5850 ;
      RECT 685.6000 319.5850 690.7500 322.5850 ;
      RECT 677.4500 319.5850 682.6000 322.5850 ;
      RECT 669.3000 319.5850 674.4500 322.5850 ;
      RECT 661.1500 319.5850 666.3000 322.5850 ;
      RECT 653.0000 319.5850 658.1500 322.5850 ;
      RECT 644.8500 319.5850 650.0000 322.5850 ;
      RECT 636.7000 319.5850 641.8500 322.5850 ;
      RECT 628.5500 319.5850 633.7000 322.5850 ;
      RECT 620.4000 319.5850 625.5500 322.5850 ;
      RECT 612.2500 319.5850 617.4000 322.5850 ;
      RECT 604.1000 319.5850 609.2500 322.5850 ;
      RECT 595.9500 319.5850 601.1000 322.5850 ;
      RECT 587.8000 319.5850 592.9500 322.5850 ;
      RECT 579.6500 319.5850 584.8000 322.5850 ;
      RECT 571.5000 319.5850 576.6500 322.5850 ;
      RECT 563.3500 319.5850 568.5000 322.5850 ;
      RECT 555.2000 319.5850 560.3500 322.5850 ;
      RECT 547.0500 319.5850 552.2000 322.5850 ;
      RECT 538.9000 319.5850 544.0500 322.5850 ;
      RECT 530.7500 319.5850 535.9000 322.5850 ;
      RECT 522.6000 319.5850 527.7500 322.5850 ;
      RECT 514.4500 319.5850 519.6000 322.5850 ;
      RECT 506.3000 319.5850 511.4500 322.5850 ;
      RECT 498.1500 319.5850 503.3000 322.5850 ;
      RECT 490.0000 319.5850 495.1500 322.5850 ;
      RECT 481.8500 319.5850 487.0000 322.5850 ;
      RECT 473.7000 319.5850 478.8500 322.5850 ;
      RECT 465.5500 319.5850 470.7000 322.5850 ;
      RECT 457.4000 319.5850 462.5500 322.5850 ;
      RECT 449.2500 319.5850 454.4000 322.5850 ;
      RECT 441.1000 319.5850 446.2500 322.5850 ;
      RECT 432.9500 319.5850 438.1000 322.5850 ;
      RECT 424.8000 319.5850 429.9500 322.5850 ;
      RECT 416.6500 319.5850 421.8000 322.5850 ;
      RECT 396.5000 319.5850 413.6500 322.5850 ;
      RECT 346.5000 319.5850 393.5000 322.5850 ;
      RECT 326.4650 319.5850 343.5000 322.5850 ;
      RECT 317.9500 319.5850 323.4650 322.5850 ;
      RECT 309.4350 319.5850 314.9500 322.5850 ;
      RECT 300.9200 319.5850 306.4350 322.5850 ;
      RECT 292.4050 319.5850 297.9200 322.5850 ;
      RECT 283.8900 319.5850 289.4050 322.5850 ;
      RECT 275.3750 319.5850 280.8900 322.5850 ;
      RECT 266.8600 319.5850 272.3750 322.5850 ;
      RECT 258.3450 319.5850 263.8600 322.5850 ;
      RECT 249.8300 319.5850 255.3450 322.5850 ;
      RECT 241.3150 319.5850 246.8300 322.5850 ;
      RECT 232.8000 319.5850 238.3150 322.5850 ;
      RECT 224.2850 319.5850 229.8000 322.5850 ;
      RECT 215.7700 319.5850 221.2850 322.5850 ;
      RECT 207.2550 319.5850 212.7700 322.5850 ;
      RECT 198.7400 319.5850 204.2550 322.5850 ;
      RECT 190.2250 319.5850 195.7400 322.5850 ;
      RECT 181.7100 319.5850 187.2250 322.5850 ;
      RECT 173.1950 319.5850 178.7100 322.5850 ;
      RECT 164.6800 319.5850 170.1950 322.5850 ;
      RECT 156.1650 319.5850 161.6800 322.5850 ;
      RECT 147.6500 319.5850 153.1650 322.5850 ;
      RECT 139.1350 319.5850 144.6500 322.5850 ;
      RECT 130.6200 319.5850 136.1350 322.5850 ;
      RECT 122.1050 319.5850 127.6200 322.5850 ;
      RECT 113.5900 319.5850 119.1050 322.5850 ;
      RECT 105.0750 319.5850 110.5900 322.5850 ;
      RECT 96.5600 319.5850 102.0750 322.5850 ;
      RECT 88.0450 319.5850 93.5600 322.5850 ;
      RECT 79.5300 319.5850 85.0450 322.5850 ;
      RECT 71.0150 319.5850 76.5300 322.5850 ;
      RECT 62.5000 319.5850 68.0150 322.5850 ;
      RECT 46.5000 319.5850 59.5000 322.5850 ;
      RECT 8.5000 319.5850 43.5000 322.5850 ;
      RECT 0.0000 319.5850 5.5000 322.5850 ;
      RECT 0.0000 318.1000 1120.0000 319.5850 ;
      RECT 1116.6000 317.5850 1120.0000 318.1000 ;
      RECT 0.0000 315.4900 1113.6000 318.1000 ;
      RECT 1118.5000 314.5850 1120.0000 317.5850 ;
      RECT 1114.5000 312.4900 1120.0000 314.5850 ;
      RECT 1076.5000 312.4900 1111.5000 315.4900 ;
      RECT 1060.5000 312.4900 1073.5000 315.4900 ;
      RECT 1052.3500 312.4900 1057.5000 315.4900 ;
      RECT 1044.2000 312.4900 1049.3500 315.4900 ;
      RECT 1036.0500 312.4900 1041.2000 315.4900 ;
      RECT 1027.9000 312.4900 1033.0500 315.4900 ;
      RECT 1019.7500 312.4900 1024.9000 315.4900 ;
      RECT 1011.6000 312.4900 1016.7500 315.4900 ;
      RECT 1003.4500 312.4900 1008.6000 315.4900 ;
      RECT 995.3000 312.4900 1000.4500 315.4900 ;
      RECT 987.1500 312.4900 992.3000 315.4900 ;
      RECT 979.0000 312.4900 984.1500 315.4900 ;
      RECT 970.8500 312.4900 976.0000 315.4900 ;
      RECT 962.7000 312.4900 967.8500 315.4900 ;
      RECT 954.5500 312.4900 959.7000 315.4900 ;
      RECT 946.4000 312.4900 951.5500 315.4900 ;
      RECT 938.2500 312.4900 943.4000 315.4900 ;
      RECT 930.1000 312.4900 935.2500 315.4900 ;
      RECT 921.9500 312.4900 927.1000 315.4900 ;
      RECT 913.8000 312.4900 918.9500 315.4900 ;
      RECT 905.6500 312.4900 910.8000 315.4900 ;
      RECT 897.5000 312.4900 902.6500 315.4900 ;
      RECT 889.3500 312.4900 894.5000 315.4900 ;
      RECT 881.2000 312.4900 886.3500 315.4900 ;
      RECT 873.0500 312.4900 878.2000 315.4900 ;
      RECT 864.9000 312.4900 870.0500 315.4900 ;
      RECT 856.7500 312.4900 861.9000 315.4900 ;
      RECT 848.6000 312.4900 853.7500 315.4900 ;
      RECT 840.4500 312.4900 845.6000 315.4900 ;
      RECT 832.3000 312.4900 837.4500 315.4900 ;
      RECT 824.1500 312.4900 829.3000 315.4900 ;
      RECT 816.0000 312.4900 821.1500 315.4900 ;
      RECT 807.8500 312.4900 813.0000 315.4900 ;
      RECT 799.7000 312.4900 804.8500 315.4900 ;
      RECT 791.5500 312.4900 796.7000 315.4900 ;
      RECT 783.4000 312.4900 788.5500 315.4900 ;
      RECT 775.2500 312.4900 780.4000 315.4900 ;
      RECT 767.1000 312.4900 772.2500 315.4900 ;
      RECT 758.9500 312.4900 764.1000 315.4900 ;
      RECT 750.8000 312.4900 755.9500 315.4900 ;
      RECT 742.6500 312.4900 747.8000 315.4900 ;
      RECT 734.5000 312.4900 739.6500 315.4900 ;
      RECT 726.3500 312.4900 731.5000 315.4900 ;
      RECT 718.2000 312.4900 723.3500 315.4900 ;
      RECT 710.0500 312.4900 715.2000 315.4900 ;
      RECT 701.9000 312.4900 707.0500 315.4900 ;
      RECT 693.7500 312.4900 698.9000 315.4900 ;
      RECT 685.6000 312.4900 690.7500 315.4900 ;
      RECT 677.4500 312.4900 682.6000 315.4900 ;
      RECT 669.3000 312.4900 674.4500 315.4900 ;
      RECT 661.1500 312.4900 666.3000 315.4900 ;
      RECT 653.0000 312.4900 658.1500 315.4900 ;
      RECT 644.8500 312.4900 650.0000 315.4900 ;
      RECT 636.7000 312.4900 641.8500 315.4900 ;
      RECT 628.5500 312.4900 633.7000 315.4900 ;
      RECT 620.4000 312.4900 625.5500 315.4900 ;
      RECT 612.2500 312.4900 617.4000 315.4900 ;
      RECT 604.1000 312.4900 609.2500 315.4900 ;
      RECT 595.9500 312.4900 601.1000 315.4900 ;
      RECT 587.8000 312.4900 592.9500 315.4900 ;
      RECT 579.6500 312.4900 584.8000 315.4900 ;
      RECT 571.5000 312.4900 576.6500 315.4900 ;
      RECT 563.3500 312.4900 568.5000 315.4900 ;
      RECT 555.2000 312.4900 560.3500 315.4900 ;
      RECT 547.0500 312.4900 552.2000 315.4900 ;
      RECT 538.9000 312.4900 544.0500 315.4900 ;
      RECT 530.7500 312.4900 535.9000 315.4900 ;
      RECT 522.6000 312.4900 527.7500 315.4900 ;
      RECT 514.4500 312.4900 519.6000 315.4900 ;
      RECT 506.3000 312.4900 511.4500 315.4900 ;
      RECT 498.1500 312.4900 503.3000 315.4900 ;
      RECT 490.0000 312.4900 495.1500 315.4900 ;
      RECT 481.8500 312.4900 487.0000 315.4900 ;
      RECT 473.7000 312.4900 478.8500 315.4900 ;
      RECT 465.5500 312.4900 470.7000 315.4900 ;
      RECT 457.4000 312.4900 462.5500 315.4900 ;
      RECT 449.2500 312.4900 454.4000 315.4900 ;
      RECT 441.1000 312.4900 446.2500 315.4900 ;
      RECT 432.9500 312.4900 438.1000 315.4900 ;
      RECT 424.8000 312.4900 429.9500 315.4900 ;
      RECT 416.6500 312.4900 421.8000 315.4900 ;
      RECT 396.5000 312.4900 413.6500 315.4900 ;
      RECT 346.5000 312.4900 393.5000 315.4900 ;
      RECT 326.4650 312.4900 343.5000 315.4900 ;
      RECT 317.9500 312.4900 323.4650 315.4900 ;
      RECT 309.4350 312.4900 314.9500 315.4900 ;
      RECT 300.9200 312.4900 306.4350 315.4900 ;
      RECT 292.4050 312.4900 297.9200 315.4900 ;
      RECT 283.8900 312.4900 289.4050 315.4900 ;
      RECT 275.3750 312.4900 280.8900 315.4900 ;
      RECT 266.8600 312.4900 272.3750 315.4900 ;
      RECT 258.3450 312.4900 263.8600 315.4900 ;
      RECT 249.8300 312.4900 255.3450 315.4900 ;
      RECT 241.3150 312.4900 246.8300 315.4900 ;
      RECT 232.8000 312.4900 238.3150 315.4900 ;
      RECT 224.2850 312.4900 229.8000 315.4900 ;
      RECT 215.7700 312.4900 221.2850 315.4900 ;
      RECT 207.2550 312.4900 212.7700 315.4900 ;
      RECT 198.7400 312.4900 204.2550 315.4900 ;
      RECT 190.2250 312.4900 195.7400 315.4900 ;
      RECT 181.7100 312.4900 187.2250 315.4900 ;
      RECT 173.1950 312.4900 178.7100 315.4900 ;
      RECT 164.6800 312.4900 170.1950 315.4900 ;
      RECT 156.1650 312.4900 161.6800 315.4900 ;
      RECT 147.6500 312.4900 153.1650 315.4900 ;
      RECT 139.1350 312.4900 144.6500 315.4900 ;
      RECT 130.6200 312.4900 136.1350 315.4900 ;
      RECT 122.1050 312.4900 127.6200 315.4900 ;
      RECT 113.5900 312.4900 119.1050 315.4900 ;
      RECT 105.0750 312.4900 110.5900 315.4900 ;
      RECT 96.5600 312.4900 102.0750 315.4900 ;
      RECT 88.0450 312.4900 93.5600 315.4900 ;
      RECT 79.5300 312.4900 85.0450 315.4900 ;
      RECT 71.0150 312.4900 76.5300 315.4900 ;
      RECT 62.5000 312.4900 68.0150 315.4900 ;
      RECT 46.5000 312.4900 59.5000 315.4900 ;
      RECT 8.5000 312.4900 43.5000 315.4900 ;
      RECT 0.0000 312.4900 5.5000 315.4900 ;
      RECT 0.0000 310.9000 1120.0000 312.4900 ;
      RECT 1116.6000 310.4900 1120.0000 310.9000 ;
      RECT 0.0000 308.3950 1113.6000 310.9000 ;
      RECT 1118.5000 307.4900 1120.0000 310.4900 ;
      RECT 1114.5000 305.3950 1120.0000 307.4900 ;
      RECT 1076.5000 305.3950 1111.5000 308.3950 ;
      RECT 1060.5000 305.3950 1073.5000 308.3950 ;
      RECT 1052.3500 305.3950 1057.5000 308.3950 ;
      RECT 1044.2000 305.3950 1049.3500 308.3950 ;
      RECT 1036.0500 305.3950 1041.2000 308.3950 ;
      RECT 1027.9000 305.3950 1033.0500 308.3950 ;
      RECT 1019.7500 305.3950 1024.9000 308.3950 ;
      RECT 1011.6000 305.3950 1016.7500 308.3950 ;
      RECT 1003.4500 305.3950 1008.6000 308.3950 ;
      RECT 995.3000 305.3950 1000.4500 308.3950 ;
      RECT 987.1500 305.3950 992.3000 308.3950 ;
      RECT 979.0000 305.3950 984.1500 308.3950 ;
      RECT 970.8500 305.3950 976.0000 308.3950 ;
      RECT 962.7000 305.3950 967.8500 308.3950 ;
      RECT 954.5500 305.3950 959.7000 308.3950 ;
      RECT 946.4000 305.3950 951.5500 308.3950 ;
      RECT 938.2500 305.3950 943.4000 308.3950 ;
      RECT 930.1000 305.3950 935.2500 308.3950 ;
      RECT 921.9500 305.3950 927.1000 308.3950 ;
      RECT 913.8000 305.3950 918.9500 308.3950 ;
      RECT 905.6500 305.3950 910.8000 308.3950 ;
      RECT 897.5000 305.3950 902.6500 308.3950 ;
      RECT 889.3500 305.3950 894.5000 308.3950 ;
      RECT 881.2000 305.3950 886.3500 308.3950 ;
      RECT 873.0500 305.3950 878.2000 308.3950 ;
      RECT 864.9000 305.3950 870.0500 308.3950 ;
      RECT 856.7500 305.3950 861.9000 308.3950 ;
      RECT 848.6000 305.3950 853.7500 308.3950 ;
      RECT 840.4500 305.3950 845.6000 308.3950 ;
      RECT 832.3000 305.3950 837.4500 308.3950 ;
      RECT 824.1500 305.3950 829.3000 308.3950 ;
      RECT 816.0000 305.3950 821.1500 308.3950 ;
      RECT 807.8500 305.3950 813.0000 308.3950 ;
      RECT 799.7000 305.3950 804.8500 308.3950 ;
      RECT 791.5500 305.3950 796.7000 308.3950 ;
      RECT 783.4000 305.3950 788.5500 308.3950 ;
      RECT 775.2500 305.3950 780.4000 308.3950 ;
      RECT 767.1000 305.3950 772.2500 308.3950 ;
      RECT 758.9500 305.3950 764.1000 308.3950 ;
      RECT 750.8000 305.3950 755.9500 308.3950 ;
      RECT 742.6500 305.3950 747.8000 308.3950 ;
      RECT 734.5000 305.3950 739.6500 308.3950 ;
      RECT 726.3500 305.3950 731.5000 308.3950 ;
      RECT 718.2000 305.3950 723.3500 308.3950 ;
      RECT 710.0500 305.3950 715.2000 308.3950 ;
      RECT 701.9000 305.3950 707.0500 308.3950 ;
      RECT 693.7500 305.3950 698.9000 308.3950 ;
      RECT 685.6000 305.3950 690.7500 308.3950 ;
      RECT 677.4500 305.3950 682.6000 308.3950 ;
      RECT 669.3000 305.3950 674.4500 308.3950 ;
      RECT 661.1500 305.3950 666.3000 308.3950 ;
      RECT 653.0000 305.3950 658.1500 308.3950 ;
      RECT 644.8500 305.3950 650.0000 308.3950 ;
      RECT 636.7000 305.3950 641.8500 308.3950 ;
      RECT 628.5500 305.3950 633.7000 308.3950 ;
      RECT 620.4000 305.3950 625.5500 308.3950 ;
      RECT 612.2500 305.3950 617.4000 308.3950 ;
      RECT 604.1000 305.3950 609.2500 308.3950 ;
      RECT 595.9500 305.3950 601.1000 308.3950 ;
      RECT 587.8000 305.3950 592.9500 308.3950 ;
      RECT 579.6500 305.3950 584.8000 308.3950 ;
      RECT 571.5000 305.3950 576.6500 308.3950 ;
      RECT 563.3500 305.3950 568.5000 308.3950 ;
      RECT 555.2000 305.3950 560.3500 308.3950 ;
      RECT 547.0500 305.3950 552.2000 308.3950 ;
      RECT 538.9000 305.3950 544.0500 308.3950 ;
      RECT 530.7500 305.3950 535.9000 308.3950 ;
      RECT 522.6000 305.3950 527.7500 308.3950 ;
      RECT 514.4500 305.3950 519.6000 308.3950 ;
      RECT 506.3000 305.3950 511.4500 308.3950 ;
      RECT 498.1500 305.3950 503.3000 308.3950 ;
      RECT 490.0000 305.3950 495.1500 308.3950 ;
      RECT 481.8500 305.3950 487.0000 308.3950 ;
      RECT 473.7000 305.3950 478.8500 308.3950 ;
      RECT 465.5500 305.3950 470.7000 308.3950 ;
      RECT 457.4000 305.3950 462.5500 308.3950 ;
      RECT 449.2500 305.3950 454.4000 308.3950 ;
      RECT 441.1000 305.3950 446.2500 308.3950 ;
      RECT 432.9500 305.3950 438.1000 308.3950 ;
      RECT 424.8000 305.3950 429.9500 308.3950 ;
      RECT 416.6500 305.3950 421.8000 308.3950 ;
      RECT 396.5000 305.3950 413.6500 308.3950 ;
      RECT 346.5000 305.3950 393.5000 308.3950 ;
      RECT 326.4650 305.3950 343.5000 308.3950 ;
      RECT 317.9500 305.3950 323.4650 308.3950 ;
      RECT 309.4350 305.3950 314.9500 308.3950 ;
      RECT 300.9200 305.3950 306.4350 308.3950 ;
      RECT 292.4050 305.3950 297.9200 308.3950 ;
      RECT 283.8900 305.3950 289.4050 308.3950 ;
      RECT 275.3750 305.3950 280.8900 308.3950 ;
      RECT 266.8600 305.3950 272.3750 308.3950 ;
      RECT 258.3450 305.3950 263.8600 308.3950 ;
      RECT 249.8300 305.3950 255.3450 308.3950 ;
      RECT 241.3150 305.3950 246.8300 308.3950 ;
      RECT 232.8000 305.3950 238.3150 308.3950 ;
      RECT 224.2850 305.3950 229.8000 308.3950 ;
      RECT 215.7700 305.3950 221.2850 308.3950 ;
      RECT 207.2550 305.3950 212.7700 308.3950 ;
      RECT 198.7400 305.3950 204.2550 308.3950 ;
      RECT 190.2250 305.3950 195.7400 308.3950 ;
      RECT 181.7100 305.3950 187.2250 308.3950 ;
      RECT 173.1950 305.3950 178.7100 308.3950 ;
      RECT 164.6800 305.3950 170.1950 308.3950 ;
      RECT 156.1650 305.3950 161.6800 308.3950 ;
      RECT 147.6500 305.3950 153.1650 308.3950 ;
      RECT 139.1350 305.3950 144.6500 308.3950 ;
      RECT 130.6200 305.3950 136.1350 308.3950 ;
      RECT 122.1050 305.3950 127.6200 308.3950 ;
      RECT 113.5900 305.3950 119.1050 308.3950 ;
      RECT 105.0750 305.3950 110.5900 308.3950 ;
      RECT 96.5600 305.3950 102.0750 308.3950 ;
      RECT 88.0450 305.3950 93.5600 308.3950 ;
      RECT 79.5300 305.3950 85.0450 308.3950 ;
      RECT 71.0150 305.3950 76.5300 308.3950 ;
      RECT 62.5000 305.3950 68.0150 308.3950 ;
      RECT 46.5000 305.3950 59.5000 308.3950 ;
      RECT 8.5000 305.3950 43.5000 308.3950 ;
      RECT 0.0000 305.3950 5.5000 308.3950 ;
      RECT 0.0000 303.9000 1120.0000 305.3950 ;
      RECT 1116.6000 303.3950 1120.0000 303.9000 ;
      RECT 0.0000 301.3000 1113.6000 303.9000 ;
      RECT 1118.5000 300.3950 1120.0000 303.3950 ;
      RECT 1114.5000 298.3000 1120.0000 300.3950 ;
      RECT 1076.5000 298.3000 1111.5000 301.3000 ;
      RECT 1060.5000 298.3000 1073.5000 301.3000 ;
      RECT 1052.3500 298.3000 1057.5000 301.3000 ;
      RECT 1044.2000 298.3000 1049.3500 301.3000 ;
      RECT 1036.0500 298.3000 1041.2000 301.3000 ;
      RECT 1027.9000 298.3000 1033.0500 301.3000 ;
      RECT 1019.7500 298.3000 1024.9000 301.3000 ;
      RECT 1011.6000 298.3000 1016.7500 301.3000 ;
      RECT 1003.4500 298.3000 1008.6000 301.3000 ;
      RECT 995.3000 298.3000 1000.4500 301.3000 ;
      RECT 987.1500 298.3000 992.3000 301.3000 ;
      RECT 979.0000 298.3000 984.1500 301.3000 ;
      RECT 970.8500 298.3000 976.0000 301.3000 ;
      RECT 962.7000 298.3000 967.8500 301.3000 ;
      RECT 954.5500 298.3000 959.7000 301.3000 ;
      RECT 946.4000 298.3000 951.5500 301.3000 ;
      RECT 938.2500 298.3000 943.4000 301.3000 ;
      RECT 930.1000 298.3000 935.2500 301.3000 ;
      RECT 921.9500 298.3000 927.1000 301.3000 ;
      RECT 913.8000 298.3000 918.9500 301.3000 ;
      RECT 905.6500 298.3000 910.8000 301.3000 ;
      RECT 897.5000 298.3000 902.6500 301.3000 ;
      RECT 889.3500 298.3000 894.5000 301.3000 ;
      RECT 881.2000 298.3000 886.3500 301.3000 ;
      RECT 873.0500 298.3000 878.2000 301.3000 ;
      RECT 864.9000 298.3000 870.0500 301.3000 ;
      RECT 856.7500 298.3000 861.9000 301.3000 ;
      RECT 848.6000 298.3000 853.7500 301.3000 ;
      RECT 840.4500 298.3000 845.6000 301.3000 ;
      RECT 832.3000 298.3000 837.4500 301.3000 ;
      RECT 824.1500 298.3000 829.3000 301.3000 ;
      RECT 816.0000 298.3000 821.1500 301.3000 ;
      RECT 807.8500 298.3000 813.0000 301.3000 ;
      RECT 799.7000 298.3000 804.8500 301.3000 ;
      RECT 791.5500 298.3000 796.7000 301.3000 ;
      RECT 783.4000 298.3000 788.5500 301.3000 ;
      RECT 775.2500 298.3000 780.4000 301.3000 ;
      RECT 767.1000 298.3000 772.2500 301.3000 ;
      RECT 758.9500 298.3000 764.1000 301.3000 ;
      RECT 750.8000 298.3000 755.9500 301.3000 ;
      RECT 742.6500 298.3000 747.8000 301.3000 ;
      RECT 734.5000 298.3000 739.6500 301.3000 ;
      RECT 726.3500 298.3000 731.5000 301.3000 ;
      RECT 718.2000 298.3000 723.3500 301.3000 ;
      RECT 710.0500 298.3000 715.2000 301.3000 ;
      RECT 701.9000 298.3000 707.0500 301.3000 ;
      RECT 693.7500 298.3000 698.9000 301.3000 ;
      RECT 685.6000 298.3000 690.7500 301.3000 ;
      RECT 677.4500 298.3000 682.6000 301.3000 ;
      RECT 669.3000 298.3000 674.4500 301.3000 ;
      RECT 661.1500 298.3000 666.3000 301.3000 ;
      RECT 653.0000 298.3000 658.1500 301.3000 ;
      RECT 644.8500 298.3000 650.0000 301.3000 ;
      RECT 636.7000 298.3000 641.8500 301.3000 ;
      RECT 628.5500 298.3000 633.7000 301.3000 ;
      RECT 620.4000 298.3000 625.5500 301.3000 ;
      RECT 612.2500 298.3000 617.4000 301.3000 ;
      RECT 604.1000 298.3000 609.2500 301.3000 ;
      RECT 595.9500 298.3000 601.1000 301.3000 ;
      RECT 587.8000 298.3000 592.9500 301.3000 ;
      RECT 579.6500 298.3000 584.8000 301.3000 ;
      RECT 571.5000 298.3000 576.6500 301.3000 ;
      RECT 563.3500 298.3000 568.5000 301.3000 ;
      RECT 555.2000 298.3000 560.3500 301.3000 ;
      RECT 547.0500 298.3000 552.2000 301.3000 ;
      RECT 538.9000 298.3000 544.0500 301.3000 ;
      RECT 530.7500 298.3000 535.9000 301.3000 ;
      RECT 522.6000 298.3000 527.7500 301.3000 ;
      RECT 514.4500 298.3000 519.6000 301.3000 ;
      RECT 506.3000 298.3000 511.4500 301.3000 ;
      RECT 498.1500 298.3000 503.3000 301.3000 ;
      RECT 490.0000 298.3000 495.1500 301.3000 ;
      RECT 481.8500 298.3000 487.0000 301.3000 ;
      RECT 473.7000 298.3000 478.8500 301.3000 ;
      RECT 465.5500 298.3000 470.7000 301.3000 ;
      RECT 457.4000 298.3000 462.5500 301.3000 ;
      RECT 449.2500 298.3000 454.4000 301.3000 ;
      RECT 441.1000 298.3000 446.2500 301.3000 ;
      RECT 432.9500 298.3000 438.1000 301.3000 ;
      RECT 424.8000 298.3000 429.9500 301.3000 ;
      RECT 416.6500 298.3000 421.8000 301.3000 ;
      RECT 396.5000 298.3000 413.6500 301.3000 ;
      RECT 346.5000 298.3000 393.5000 301.3000 ;
      RECT 326.4650 298.3000 343.5000 301.3000 ;
      RECT 317.9500 298.3000 323.4650 301.3000 ;
      RECT 309.4350 298.3000 314.9500 301.3000 ;
      RECT 300.9200 298.3000 306.4350 301.3000 ;
      RECT 292.4050 298.3000 297.9200 301.3000 ;
      RECT 283.8900 298.3000 289.4050 301.3000 ;
      RECT 275.3750 298.3000 280.8900 301.3000 ;
      RECT 266.8600 298.3000 272.3750 301.3000 ;
      RECT 258.3450 298.3000 263.8600 301.3000 ;
      RECT 249.8300 298.3000 255.3450 301.3000 ;
      RECT 241.3150 298.3000 246.8300 301.3000 ;
      RECT 232.8000 298.3000 238.3150 301.3000 ;
      RECT 224.2850 298.3000 229.8000 301.3000 ;
      RECT 215.7700 298.3000 221.2850 301.3000 ;
      RECT 207.2550 298.3000 212.7700 301.3000 ;
      RECT 198.7400 298.3000 204.2550 301.3000 ;
      RECT 190.2250 298.3000 195.7400 301.3000 ;
      RECT 181.7100 298.3000 187.2250 301.3000 ;
      RECT 173.1950 298.3000 178.7100 301.3000 ;
      RECT 164.6800 298.3000 170.1950 301.3000 ;
      RECT 156.1650 298.3000 161.6800 301.3000 ;
      RECT 147.6500 298.3000 153.1650 301.3000 ;
      RECT 139.1350 298.3000 144.6500 301.3000 ;
      RECT 130.6200 298.3000 136.1350 301.3000 ;
      RECT 122.1050 298.3000 127.6200 301.3000 ;
      RECT 113.5900 298.3000 119.1050 301.3000 ;
      RECT 105.0750 298.3000 110.5900 301.3000 ;
      RECT 96.5600 298.3000 102.0750 301.3000 ;
      RECT 88.0450 298.3000 93.5600 301.3000 ;
      RECT 79.5300 298.3000 85.0450 301.3000 ;
      RECT 71.0150 298.3000 76.5300 301.3000 ;
      RECT 62.5000 298.3000 68.0150 301.3000 ;
      RECT 46.5000 298.3000 59.5000 301.3000 ;
      RECT 8.5000 298.3000 43.5000 301.3000 ;
      RECT 0.0000 298.3000 5.5000 301.3000 ;
      RECT 0.0000 296.9000 1120.0000 298.3000 ;
      RECT 1116.6000 296.3000 1120.0000 296.9000 ;
      RECT 0.0000 294.2050 1113.6000 296.9000 ;
      RECT 1118.5000 293.3000 1120.0000 296.3000 ;
      RECT 1114.5000 291.2050 1120.0000 293.3000 ;
      RECT 1076.5000 291.2050 1111.5000 294.2050 ;
      RECT 1060.5000 291.2050 1073.5000 294.2050 ;
      RECT 1052.3500 291.2050 1057.5000 294.2050 ;
      RECT 1044.2000 291.2050 1049.3500 294.2050 ;
      RECT 1036.0500 291.2050 1041.2000 294.2050 ;
      RECT 1027.9000 291.2050 1033.0500 294.2050 ;
      RECT 1019.7500 291.2050 1024.9000 294.2050 ;
      RECT 1011.6000 291.2050 1016.7500 294.2050 ;
      RECT 1003.4500 291.2050 1008.6000 294.2050 ;
      RECT 995.3000 291.2050 1000.4500 294.2050 ;
      RECT 987.1500 291.2050 992.3000 294.2050 ;
      RECT 979.0000 291.2050 984.1500 294.2050 ;
      RECT 970.8500 291.2050 976.0000 294.2050 ;
      RECT 962.7000 291.2050 967.8500 294.2050 ;
      RECT 954.5500 291.2050 959.7000 294.2050 ;
      RECT 946.4000 291.2050 951.5500 294.2050 ;
      RECT 938.2500 291.2050 943.4000 294.2050 ;
      RECT 930.1000 291.2050 935.2500 294.2050 ;
      RECT 921.9500 291.2050 927.1000 294.2050 ;
      RECT 913.8000 291.2050 918.9500 294.2050 ;
      RECT 905.6500 291.2050 910.8000 294.2050 ;
      RECT 897.5000 291.2050 902.6500 294.2050 ;
      RECT 889.3500 291.2050 894.5000 294.2050 ;
      RECT 881.2000 291.2050 886.3500 294.2050 ;
      RECT 873.0500 291.2050 878.2000 294.2050 ;
      RECT 864.9000 291.2050 870.0500 294.2050 ;
      RECT 856.7500 291.2050 861.9000 294.2050 ;
      RECT 848.6000 291.2050 853.7500 294.2050 ;
      RECT 840.4500 291.2050 845.6000 294.2050 ;
      RECT 832.3000 291.2050 837.4500 294.2050 ;
      RECT 824.1500 291.2050 829.3000 294.2050 ;
      RECT 816.0000 291.2050 821.1500 294.2050 ;
      RECT 807.8500 291.2050 813.0000 294.2050 ;
      RECT 799.7000 291.2050 804.8500 294.2050 ;
      RECT 791.5500 291.2050 796.7000 294.2050 ;
      RECT 783.4000 291.2050 788.5500 294.2050 ;
      RECT 775.2500 291.2050 780.4000 294.2050 ;
      RECT 767.1000 291.2050 772.2500 294.2050 ;
      RECT 758.9500 291.2050 764.1000 294.2050 ;
      RECT 750.8000 291.2050 755.9500 294.2050 ;
      RECT 742.6500 291.2050 747.8000 294.2050 ;
      RECT 734.5000 291.2050 739.6500 294.2050 ;
      RECT 726.3500 291.2050 731.5000 294.2050 ;
      RECT 718.2000 291.2050 723.3500 294.2050 ;
      RECT 710.0500 291.2050 715.2000 294.2050 ;
      RECT 701.9000 291.2050 707.0500 294.2050 ;
      RECT 693.7500 291.2050 698.9000 294.2050 ;
      RECT 685.6000 291.2050 690.7500 294.2050 ;
      RECT 677.4500 291.2050 682.6000 294.2050 ;
      RECT 669.3000 291.2050 674.4500 294.2050 ;
      RECT 661.1500 291.2050 666.3000 294.2050 ;
      RECT 653.0000 291.2050 658.1500 294.2050 ;
      RECT 644.8500 291.2050 650.0000 294.2050 ;
      RECT 636.7000 291.2050 641.8500 294.2050 ;
      RECT 628.5500 291.2050 633.7000 294.2050 ;
      RECT 620.4000 291.2050 625.5500 294.2050 ;
      RECT 612.2500 291.2050 617.4000 294.2050 ;
      RECT 604.1000 291.2050 609.2500 294.2050 ;
      RECT 595.9500 291.2050 601.1000 294.2050 ;
      RECT 587.8000 291.2050 592.9500 294.2050 ;
      RECT 579.6500 291.2050 584.8000 294.2050 ;
      RECT 571.5000 291.2050 576.6500 294.2050 ;
      RECT 563.3500 291.2050 568.5000 294.2050 ;
      RECT 555.2000 291.2050 560.3500 294.2050 ;
      RECT 547.0500 291.2050 552.2000 294.2050 ;
      RECT 538.9000 291.2050 544.0500 294.2050 ;
      RECT 530.7500 291.2050 535.9000 294.2050 ;
      RECT 522.6000 291.2050 527.7500 294.2050 ;
      RECT 514.4500 291.2050 519.6000 294.2050 ;
      RECT 506.3000 291.2050 511.4500 294.2050 ;
      RECT 498.1500 291.2050 503.3000 294.2050 ;
      RECT 490.0000 291.2050 495.1500 294.2050 ;
      RECT 481.8500 291.2050 487.0000 294.2050 ;
      RECT 473.7000 291.2050 478.8500 294.2050 ;
      RECT 465.5500 291.2050 470.7000 294.2050 ;
      RECT 457.4000 291.2050 462.5500 294.2050 ;
      RECT 449.2500 291.2050 454.4000 294.2050 ;
      RECT 441.1000 291.2050 446.2500 294.2050 ;
      RECT 432.9500 291.2050 438.1000 294.2050 ;
      RECT 424.8000 291.2050 429.9500 294.2050 ;
      RECT 416.6500 291.2050 421.8000 294.2050 ;
      RECT 396.5000 291.2050 413.6500 294.2050 ;
      RECT 346.5000 291.2050 393.5000 294.2050 ;
      RECT 326.4650 291.2050 343.5000 294.2050 ;
      RECT 317.9500 291.2050 323.4650 294.2050 ;
      RECT 309.4350 291.2050 314.9500 294.2050 ;
      RECT 300.9200 291.2050 306.4350 294.2050 ;
      RECT 292.4050 291.2050 297.9200 294.2050 ;
      RECT 283.8900 291.2050 289.4050 294.2050 ;
      RECT 275.3750 291.2050 280.8900 294.2050 ;
      RECT 266.8600 291.2050 272.3750 294.2050 ;
      RECT 258.3450 291.2050 263.8600 294.2050 ;
      RECT 249.8300 291.2050 255.3450 294.2050 ;
      RECT 241.3150 291.2050 246.8300 294.2050 ;
      RECT 232.8000 291.2050 238.3150 294.2050 ;
      RECT 224.2850 291.2050 229.8000 294.2050 ;
      RECT 215.7700 291.2050 221.2850 294.2050 ;
      RECT 207.2550 291.2050 212.7700 294.2050 ;
      RECT 198.7400 291.2050 204.2550 294.2050 ;
      RECT 190.2250 291.2050 195.7400 294.2050 ;
      RECT 181.7100 291.2050 187.2250 294.2050 ;
      RECT 173.1950 291.2050 178.7100 294.2050 ;
      RECT 164.6800 291.2050 170.1950 294.2050 ;
      RECT 156.1650 291.2050 161.6800 294.2050 ;
      RECT 147.6500 291.2050 153.1650 294.2050 ;
      RECT 139.1350 291.2050 144.6500 294.2050 ;
      RECT 130.6200 291.2050 136.1350 294.2050 ;
      RECT 122.1050 291.2050 127.6200 294.2050 ;
      RECT 113.5900 291.2050 119.1050 294.2050 ;
      RECT 105.0750 291.2050 110.5900 294.2050 ;
      RECT 96.5600 291.2050 102.0750 294.2050 ;
      RECT 88.0450 291.2050 93.5600 294.2050 ;
      RECT 79.5300 291.2050 85.0450 294.2050 ;
      RECT 71.0150 291.2050 76.5300 294.2050 ;
      RECT 62.5000 291.2050 68.0150 294.2050 ;
      RECT 46.5000 291.2050 59.5000 294.2050 ;
      RECT 8.5000 291.2050 43.5000 294.2050 ;
      RECT 0.0000 291.2050 5.5000 294.2050 ;
      RECT 0.0000 289.7000 1120.0000 291.2050 ;
      RECT 1116.6000 289.2050 1120.0000 289.7000 ;
      RECT 0.0000 287.1100 1113.6000 289.7000 ;
      RECT 1118.5000 286.2050 1120.0000 289.2050 ;
      RECT 1114.5000 284.1100 1120.0000 286.2050 ;
      RECT 1076.5000 284.1100 1111.5000 287.1100 ;
      RECT 1060.5000 284.1100 1073.5000 287.1100 ;
      RECT 1052.3500 284.1100 1057.5000 287.1100 ;
      RECT 1044.2000 284.1100 1049.3500 287.1100 ;
      RECT 1036.0500 284.1100 1041.2000 287.1100 ;
      RECT 1027.9000 284.1100 1033.0500 287.1100 ;
      RECT 1019.7500 284.1100 1024.9000 287.1100 ;
      RECT 1011.6000 284.1100 1016.7500 287.1100 ;
      RECT 1003.4500 284.1100 1008.6000 287.1100 ;
      RECT 995.3000 284.1100 1000.4500 287.1100 ;
      RECT 987.1500 284.1100 992.3000 287.1100 ;
      RECT 979.0000 284.1100 984.1500 287.1100 ;
      RECT 970.8500 284.1100 976.0000 287.1100 ;
      RECT 962.7000 284.1100 967.8500 287.1100 ;
      RECT 954.5500 284.1100 959.7000 287.1100 ;
      RECT 946.4000 284.1100 951.5500 287.1100 ;
      RECT 938.2500 284.1100 943.4000 287.1100 ;
      RECT 930.1000 284.1100 935.2500 287.1100 ;
      RECT 921.9500 284.1100 927.1000 287.1100 ;
      RECT 913.8000 284.1100 918.9500 287.1100 ;
      RECT 905.6500 284.1100 910.8000 287.1100 ;
      RECT 897.5000 284.1100 902.6500 287.1100 ;
      RECT 889.3500 284.1100 894.5000 287.1100 ;
      RECT 881.2000 284.1100 886.3500 287.1100 ;
      RECT 873.0500 284.1100 878.2000 287.1100 ;
      RECT 864.9000 284.1100 870.0500 287.1100 ;
      RECT 856.7500 284.1100 861.9000 287.1100 ;
      RECT 848.6000 284.1100 853.7500 287.1100 ;
      RECT 840.4500 284.1100 845.6000 287.1100 ;
      RECT 832.3000 284.1100 837.4500 287.1100 ;
      RECT 824.1500 284.1100 829.3000 287.1100 ;
      RECT 816.0000 284.1100 821.1500 287.1100 ;
      RECT 807.8500 284.1100 813.0000 287.1100 ;
      RECT 799.7000 284.1100 804.8500 287.1100 ;
      RECT 791.5500 284.1100 796.7000 287.1100 ;
      RECT 783.4000 284.1100 788.5500 287.1100 ;
      RECT 775.2500 284.1100 780.4000 287.1100 ;
      RECT 767.1000 284.1100 772.2500 287.1100 ;
      RECT 758.9500 284.1100 764.1000 287.1100 ;
      RECT 750.8000 284.1100 755.9500 287.1100 ;
      RECT 742.6500 284.1100 747.8000 287.1100 ;
      RECT 734.5000 284.1100 739.6500 287.1100 ;
      RECT 726.3500 284.1100 731.5000 287.1100 ;
      RECT 718.2000 284.1100 723.3500 287.1100 ;
      RECT 710.0500 284.1100 715.2000 287.1100 ;
      RECT 701.9000 284.1100 707.0500 287.1100 ;
      RECT 693.7500 284.1100 698.9000 287.1100 ;
      RECT 685.6000 284.1100 690.7500 287.1100 ;
      RECT 677.4500 284.1100 682.6000 287.1100 ;
      RECT 669.3000 284.1100 674.4500 287.1100 ;
      RECT 661.1500 284.1100 666.3000 287.1100 ;
      RECT 653.0000 284.1100 658.1500 287.1100 ;
      RECT 644.8500 284.1100 650.0000 287.1100 ;
      RECT 636.7000 284.1100 641.8500 287.1100 ;
      RECT 628.5500 284.1100 633.7000 287.1100 ;
      RECT 620.4000 284.1100 625.5500 287.1100 ;
      RECT 612.2500 284.1100 617.4000 287.1100 ;
      RECT 604.1000 284.1100 609.2500 287.1100 ;
      RECT 595.9500 284.1100 601.1000 287.1100 ;
      RECT 587.8000 284.1100 592.9500 287.1100 ;
      RECT 579.6500 284.1100 584.8000 287.1100 ;
      RECT 571.5000 284.1100 576.6500 287.1100 ;
      RECT 563.3500 284.1100 568.5000 287.1100 ;
      RECT 555.2000 284.1100 560.3500 287.1100 ;
      RECT 547.0500 284.1100 552.2000 287.1100 ;
      RECT 538.9000 284.1100 544.0500 287.1100 ;
      RECT 530.7500 284.1100 535.9000 287.1100 ;
      RECT 522.6000 284.1100 527.7500 287.1100 ;
      RECT 514.4500 284.1100 519.6000 287.1100 ;
      RECT 506.3000 284.1100 511.4500 287.1100 ;
      RECT 498.1500 284.1100 503.3000 287.1100 ;
      RECT 490.0000 284.1100 495.1500 287.1100 ;
      RECT 481.8500 284.1100 487.0000 287.1100 ;
      RECT 473.7000 284.1100 478.8500 287.1100 ;
      RECT 465.5500 284.1100 470.7000 287.1100 ;
      RECT 457.4000 284.1100 462.5500 287.1100 ;
      RECT 449.2500 284.1100 454.4000 287.1100 ;
      RECT 441.1000 284.1100 446.2500 287.1100 ;
      RECT 432.9500 284.1100 438.1000 287.1100 ;
      RECT 424.8000 284.1100 429.9500 287.1100 ;
      RECT 416.6500 284.1100 421.8000 287.1100 ;
      RECT 396.5000 284.1100 413.6500 287.1100 ;
      RECT 346.5000 284.1100 393.5000 287.1100 ;
      RECT 326.4650 284.1100 343.5000 287.1100 ;
      RECT 317.9500 284.1100 323.4650 287.1100 ;
      RECT 309.4350 284.1100 314.9500 287.1100 ;
      RECT 300.9200 284.1100 306.4350 287.1100 ;
      RECT 292.4050 284.1100 297.9200 287.1100 ;
      RECT 283.8900 284.1100 289.4050 287.1100 ;
      RECT 275.3750 284.1100 280.8900 287.1100 ;
      RECT 266.8600 284.1100 272.3750 287.1100 ;
      RECT 258.3450 284.1100 263.8600 287.1100 ;
      RECT 249.8300 284.1100 255.3450 287.1100 ;
      RECT 241.3150 284.1100 246.8300 287.1100 ;
      RECT 232.8000 284.1100 238.3150 287.1100 ;
      RECT 224.2850 284.1100 229.8000 287.1100 ;
      RECT 215.7700 284.1100 221.2850 287.1100 ;
      RECT 207.2550 284.1100 212.7700 287.1100 ;
      RECT 198.7400 284.1100 204.2550 287.1100 ;
      RECT 190.2250 284.1100 195.7400 287.1100 ;
      RECT 181.7100 284.1100 187.2250 287.1100 ;
      RECT 173.1950 284.1100 178.7100 287.1100 ;
      RECT 164.6800 284.1100 170.1950 287.1100 ;
      RECT 156.1650 284.1100 161.6800 287.1100 ;
      RECT 147.6500 284.1100 153.1650 287.1100 ;
      RECT 139.1350 284.1100 144.6500 287.1100 ;
      RECT 130.6200 284.1100 136.1350 287.1100 ;
      RECT 122.1050 284.1100 127.6200 287.1100 ;
      RECT 113.5900 284.1100 119.1050 287.1100 ;
      RECT 105.0750 284.1100 110.5900 287.1100 ;
      RECT 96.5600 284.1100 102.0750 287.1100 ;
      RECT 88.0450 284.1100 93.5600 287.1100 ;
      RECT 79.5300 284.1100 85.0450 287.1100 ;
      RECT 71.0150 284.1100 76.5300 287.1100 ;
      RECT 62.5000 284.1100 68.0150 287.1100 ;
      RECT 46.5000 284.1100 59.5000 287.1100 ;
      RECT 8.5000 284.1100 43.5000 287.1100 ;
      RECT 0.0000 284.1100 5.5000 287.1100 ;
      RECT 0.0000 283.3000 1120.0000 284.1100 ;
      RECT 1116.6000 282.1100 1120.0000 283.3000 ;
      RECT 0.0000 280.0150 1113.6000 283.3000 ;
      RECT 1118.5000 279.1100 1120.0000 282.1100 ;
      RECT 1114.5000 277.0150 1120.0000 279.1100 ;
      RECT 1076.5000 277.0150 1111.5000 280.0150 ;
      RECT 1060.5000 277.0150 1073.5000 280.0150 ;
      RECT 1052.3500 277.0150 1057.5000 280.0150 ;
      RECT 1044.2000 277.0150 1049.3500 280.0150 ;
      RECT 1036.0500 277.0150 1041.2000 280.0150 ;
      RECT 1027.9000 277.0150 1033.0500 280.0150 ;
      RECT 1019.7500 277.0150 1024.9000 280.0150 ;
      RECT 1011.6000 277.0150 1016.7500 280.0150 ;
      RECT 1003.4500 277.0150 1008.6000 280.0150 ;
      RECT 995.3000 277.0150 1000.4500 280.0150 ;
      RECT 987.1500 277.0150 992.3000 280.0150 ;
      RECT 979.0000 277.0150 984.1500 280.0150 ;
      RECT 970.8500 277.0150 976.0000 280.0150 ;
      RECT 962.7000 277.0150 967.8500 280.0150 ;
      RECT 954.5500 277.0150 959.7000 280.0150 ;
      RECT 946.4000 277.0150 951.5500 280.0150 ;
      RECT 938.2500 277.0150 943.4000 280.0150 ;
      RECT 930.1000 277.0150 935.2500 280.0150 ;
      RECT 921.9500 277.0150 927.1000 280.0150 ;
      RECT 913.8000 277.0150 918.9500 280.0150 ;
      RECT 905.6500 277.0150 910.8000 280.0150 ;
      RECT 897.5000 277.0150 902.6500 280.0150 ;
      RECT 889.3500 277.0150 894.5000 280.0150 ;
      RECT 881.2000 277.0150 886.3500 280.0150 ;
      RECT 873.0500 277.0150 878.2000 280.0150 ;
      RECT 864.9000 277.0150 870.0500 280.0150 ;
      RECT 856.7500 277.0150 861.9000 280.0150 ;
      RECT 848.6000 277.0150 853.7500 280.0150 ;
      RECT 840.4500 277.0150 845.6000 280.0150 ;
      RECT 832.3000 277.0150 837.4500 280.0150 ;
      RECT 824.1500 277.0150 829.3000 280.0150 ;
      RECT 816.0000 277.0150 821.1500 280.0150 ;
      RECT 807.8500 277.0150 813.0000 280.0150 ;
      RECT 799.7000 277.0150 804.8500 280.0150 ;
      RECT 791.5500 277.0150 796.7000 280.0150 ;
      RECT 783.4000 277.0150 788.5500 280.0150 ;
      RECT 775.2500 277.0150 780.4000 280.0150 ;
      RECT 767.1000 277.0150 772.2500 280.0150 ;
      RECT 758.9500 277.0150 764.1000 280.0150 ;
      RECT 750.8000 277.0150 755.9500 280.0150 ;
      RECT 742.6500 277.0150 747.8000 280.0150 ;
      RECT 734.5000 277.0150 739.6500 280.0150 ;
      RECT 726.3500 277.0150 731.5000 280.0150 ;
      RECT 718.2000 277.0150 723.3500 280.0150 ;
      RECT 710.0500 277.0150 715.2000 280.0150 ;
      RECT 701.9000 277.0150 707.0500 280.0150 ;
      RECT 693.7500 277.0150 698.9000 280.0150 ;
      RECT 685.6000 277.0150 690.7500 280.0150 ;
      RECT 677.4500 277.0150 682.6000 280.0150 ;
      RECT 669.3000 277.0150 674.4500 280.0150 ;
      RECT 661.1500 277.0150 666.3000 280.0150 ;
      RECT 653.0000 277.0150 658.1500 280.0150 ;
      RECT 644.8500 277.0150 650.0000 280.0150 ;
      RECT 636.7000 277.0150 641.8500 280.0150 ;
      RECT 628.5500 277.0150 633.7000 280.0150 ;
      RECT 620.4000 277.0150 625.5500 280.0150 ;
      RECT 612.2500 277.0150 617.4000 280.0150 ;
      RECT 604.1000 277.0150 609.2500 280.0150 ;
      RECT 595.9500 277.0150 601.1000 280.0150 ;
      RECT 587.8000 277.0150 592.9500 280.0150 ;
      RECT 579.6500 277.0150 584.8000 280.0150 ;
      RECT 571.5000 277.0150 576.6500 280.0150 ;
      RECT 563.3500 277.0150 568.5000 280.0150 ;
      RECT 555.2000 277.0150 560.3500 280.0150 ;
      RECT 547.0500 277.0150 552.2000 280.0150 ;
      RECT 538.9000 277.0150 544.0500 280.0150 ;
      RECT 530.7500 277.0150 535.9000 280.0150 ;
      RECT 522.6000 277.0150 527.7500 280.0150 ;
      RECT 514.4500 277.0150 519.6000 280.0150 ;
      RECT 506.3000 277.0150 511.4500 280.0150 ;
      RECT 498.1500 277.0150 503.3000 280.0150 ;
      RECT 490.0000 277.0150 495.1500 280.0150 ;
      RECT 481.8500 277.0150 487.0000 280.0150 ;
      RECT 473.7000 277.0150 478.8500 280.0150 ;
      RECT 465.5500 277.0150 470.7000 280.0150 ;
      RECT 457.4000 277.0150 462.5500 280.0150 ;
      RECT 449.2500 277.0150 454.4000 280.0150 ;
      RECT 441.1000 277.0150 446.2500 280.0150 ;
      RECT 432.9500 277.0150 438.1000 280.0150 ;
      RECT 424.8000 277.0150 429.9500 280.0150 ;
      RECT 416.6500 277.0150 421.8000 280.0150 ;
      RECT 396.5000 277.0150 413.6500 280.0150 ;
      RECT 346.5000 277.0150 393.5000 280.0150 ;
      RECT 326.4650 277.0150 343.5000 280.0150 ;
      RECT 317.9500 277.0150 323.4650 280.0150 ;
      RECT 309.4350 277.0150 314.9500 280.0150 ;
      RECT 300.9200 277.0150 306.4350 280.0150 ;
      RECT 292.4050 277.0150 297.9200 280.0150 ;
      RECT 283.8900 277.0150 289.4050 280.0150 ;
      RECT 275.3750 277.0150 280.8900 280.0150 ;
      RECT 266.8600 277.0150 272.3750 280.0150 ;
      RECT 258.3450 277.0150 263.8600 280.0150 ;
      RECT 249.8300 277.0150 255.3450 280.0150 ;
      RECT 241.3150 277.0150 246.8300 280.0150 ;
      RECT 232.8000 277.0150 238.3150 280.0150 ;
      RECT 224.2850 277.0150 229.8000 280.0150 ;
      RECT 215.7700 277.0150 221.2850 280.0150 ;
      RECT 207.2550 277.0150 212.7700 280.0150 ;
      RECT 198.7400 277.0150 204.2550 280.0150 ;
      RECT 190.2250 277.0150 195.7400 280.0150 ;
      RECT 181.7100 277.0150 187.2250 280.0150 ;
      RECT 173.1950 277.0150 178.7100 280.0150 ;
      RECT 164.6800 277.0150 170.1950 280.0150 ;
      RECT 156.1650 277.0150 161.6800 280.0150 ;
      RECT 147.6500 277.0150 153.1650 280.0150 ;
      RECT 139.1350 277.0150 144.6500 280.0150 ;
      RECT 130.6200 277.0150 136.1350 280.0150 ;
      RECT 122.1050 277.0150 127.6200 280.0150 ;
      RECT 113.5900 277.0150 119.1050 280.0150 ;
      RECT 105.0750 277.0150 110.5900 280.0150 ;
      RECT 96.5600 277.0150 102.0750 280.0150 ;
      RECT 88.0450 277.0150 93.5600 280.0150 ;
      RECT 79.5300 277.0150 85.0450 280.0150 ;
      RECT 71.0150 277.0150 76.5300 280.0150 ;
      RECT 62.5000 277.0150 68.0150 280.0150 ;
      RECT 46.5000 277.0150 59.5000 280.0150 ;
      RECT 8.5000 277.0150 43.5000 280.0150 ;
      RECT 0.0000 277.0150 5.5000 280.0150 ;
      RECT 0.0000 276.1000 1120.0000 277.0150 ;
      RECT 1116.6000 275.0150 1120.0000 276.1000 ;
      RECT 0.0000 272.9200 1113.6000 276.1000 ;
      RECT 1118.5000 272.0150 1120.0000 275.0150 ;
      RECT 1114.5000 269.9200 1120.0000 272.0150 ;
      RECT 1076.5000 269.9200 1111.5000 272.9200 ;
      RECT 1060.5000 269.9200 1073.5000 272.9200 ;
      RECT 1052.3500 269.9200 1057.5000 272.9200 ;
      RECT 1044.2000 269.9200 1049.3500 272.9200 ;
      RECT 1036.0500 269.9200 1041.2000 272.9200 ;
      RECT 1027.9000 269.9200 1033.0500 272.9200 ;
      RECT 1019.7500 269.9200 1024.9000 272.9200 ;
      RECT 1011.6000 269.9200 1016.7500 272.9200 ;
      RECT 1003.4500 269.9200 1008.6000 272.9200 ;
      RECT 995.3000 269.9200 1000.4500 272.9200 ;
      RECT 987.1500 269.9200 992.3000 272.9200 ;
      RECT 979.0000 269.9200 984.1500 272.9200 ;
      RECT 970.8500 269.9200 976.0000 272.9200 ;
      RECT 962.7000 269.9200 967.8500 272.9200 ;
      RECT 954.5500 269.9200 959.7000 272.9200 ;
      RECT 946.4000 269.9200 951.5500 272.9200 ;
      RECT 938.2500 269.9200 943.4000 272.9200 ;
      RECT 930.1000 269.9200 935.2500 272.9200 ;
      RECT 921.9500 269.9200 927.1000 272.9200 ;
      RECT 913.8000 269.9200 918.9500 272.9200 ;
      RECT 905.6500 269.9200 910.8000 272.9200 ;
      RECT 897.5000 269.9200 902.6500 272.9200 ;
      RECT 889.3500 269.9200 894.5000 272.9200 ;
      RECT 881.2000 269.9200 886.3500 272.9200 ;
      RECT 873.0500 269.9200 878.2000 272.9200 ;
      RECT 864.9000 269.9200 870.0500 272.9200 ;
      RECT 856.7500 269.9200 861.9000 272.9200 ;
      RECT 848.6000 269.9200 853.7500 272.9200 ;
      RECT 840.4500 269.9200 845.6000 272.9200 ;
      RECT 832.3000 269.9200 837.4500 272.9200 ;
      RECT 824.1500 269.9200 829.3000 272.9200 ;
      RECT 816.0000 269.9200 821.1500 272.9200 ;
      RECT 807.8500 269.9200 813.0000 272.9200 ;
      RECT 799.7000 269.9200 804.8500 272.9200 ;
      RECT 791.5500 269.9200 796.7000 272.9200 ;
      RECT 783.4000 269.9200 788.5500 272.9200 ;
      RECT 775.2500 269.9200 780.4000 272.9200 ;
      RECT 767.1000 269.9200 772.2500 272.9200 ;
      RECT 758.9500 269.9200 764.1000 272.9200 ;
      RECT 750.8000 269.9200 755.9500 272.9200 ;
      RECT 742.6500 269.9200 747.8000 272.9200 ;
      RECT 734.5000 269.9200 739.6500 272.9200 ;
      RECT 726.3500 269.9200 731.5000 272.9200 ;
      RECT 718.2000 269.9200 723.3500 272.9200 ;
      RECT 710.0500 269.9200 715.2000 272.9200 ;
      RECT 701.9000 269.9200 707.0500 272.9200 ;
      RECT 693.7500 269.9200 698.9000 272.9200 ;
      RECT 685.6000 269.9200 690.7500 272.9200 ;
      RECT 677.4500 269.9200 682.6000 272.9200 ;
      RECT 669.3000 269.9200 674.4500 272.9200 ;
      RECT 661.1500 269.9200 666.3000 272.9200 ;
      RECT 653.0000 269.9200 658.1500 272.9200 ;
      RECT 644.8500 269.9200 650.0000 272.9200 ;
      RECT 636.7000 269.9200 641.8500 272.9200 ;
      RECT 628.5500 269.9200 633.7000 272.9200 ;
      RECT 620.4000 269.9200 625.5500 272.9200 ;
      RECT 612.2500 269.9200 617.4000 272.9200 ;
      RECT 604.1000 269.9200 609.2500 272.9200 ;
      RECT 595.9500 269.9200 601.1000 272.9200 ;
      RECT 587.8000 269.9200 592.9500 272.9200 ;
      RECT 579.6500 269.9200 584.8000 272.9200 ;
      RECT 571.5000 269.9200 576.6500 272.9200 ;
      RECT 563.3500 269.9200 568.5000 272.9200 ;
      RECT 555.2000 269.9200 560.3500 272.9200 ;
      RECT 547.0500 269.9200 552.2000 272.9200 ;
      RECT 538.9000 269.9200 544.0500 272.9200 ;
      RECT 530.7500 269.9200 535.9000 272.9200 ;
      RECT 522.6000 269.9200 527.7500 272.9200 ;
      RECT 514.4500 269.9200 519.6000 272.9200 ;
      RECT 506.3000 269.9200 511.4500 272.9200 ;
      RECT 498.1500 269.9200 503.3000 272.9200 ;
      RECT 490.0000 269.9200 495.1500 272.9200 ;
      RECT 481.8500 269.9200 487.0000 272.9200 ;
      RECT 473.7000 269.9200 478.8500 272.9200 ;
      RECT 465.5500 269.9200 470.7000 272.9200 ;
      RECT 457.4000 269.9200 462.5500 272.9200 ;
      RECT 449.2500 269.9200 454.4000 272.9200 ;
      RECT 441.1000 269.9200 446.2500 272.9200 ;
      RECT 432.9500 269.9200 438.1000 272.9200 ;
      RECT 424.8000 269.9200 429.9500 272.9200 ;
      RECT 416.6500 269.9200 421.8000 272.9200 ;
      RECT 396.5000 269.9200 413.6500 272.9200 ;
      RECT 346.5000 269.9200 393.5000 272.9200 ;
      RECT 326.4650 269.9200 343.5000 272.9200 ;
      RECT 317.9500 269.9200 323.4650 272.9200 ;
      RECT 309.4350 269.9200 314.9500 272.9200 ;
      RECT 300.9200 269.9200 306.4350 272.9200 ;
      RECT 292.4050 269.9200 297.9200 272.9200 ;
      RECT 283.8900 269.9200 289.4050 272.9200 ;
      RECT 275.3750 269.9200 280.8900 272.9200 ;
      RECT 266.8600 269.9200 272.3750 272.9200 ;
      RECT 258.3450 269.9200 263.8600 272.9200 ;
      RECT 249.8300 269.9200 255.3450 272.9200 ;
      RECT 241.3150 269.9200 246.8300 272.9200 ;
      RECT 232.8000 269.9200 238.3150 272.9200 ;
      RECT 224.2850 269.9200 229.8000 272.9200 ;
      RECT 215.7700 269.9200 221.2850 272.9200 ;
      RECT 207.2550 269.9200 212.7700 272.9200 ;
      RECT 198.7400 269.9200 204.2550 272.9200 ;
      RECT 190.2250 269.9200 195.7400 272.9200 ;
      RECT 181.7100 269.9200 187.2250 272.9200 ;
      RECT 173.1950 269.9200 178.7100 272.9200 ;
      RECT 164.6800 269.9200 170.1950 272.9200 ;
      RECT 156.1650 269.9200 161.6800 272.9200 ;
      RECT 147.6500 269.9200 153.1650 272.9200 ;
      RECT 139.1350 269.9200 144.6500 272.9200 ;
      RECT 130.6200 269.9200 136.1350 272.9200 ;
      RECT 122.1050 269.9200 127.6200 272.9200 ;
      RECT 113.5900 269.9200 119.1050 272.9200 ;
      RECT 105.0750 269.9200 110.5900 272.9200 ;
      RECT 96.5600 269.9200 102.0750 272.9200 ;
      RECT 88.0450 269.9200 93.5600 272.9200 ;
      RECT 79.5300 269.9200 85.0450 272.9200 ;
      RECT 71.0150 269.9200 76.5300 272.9200 ;
      RECT 62.5000 269.9200 68.0150 272.9200 ;
      RECT 46.5000 269.9200 59.5000 272.9200 ;
      RECT 8.5000 269.9200 43.5000 272.9200 ;
      RECT 0.0000 269.9200 5.5000 272.9200 ;
      RECT 0.0000 268.9000 1120.0000 269.9200 ;
      RECT 1116.6000 267.9200 1120.0000 268.9000 ;
      RECT 0.0000 265.8250 1113.6000 268.9000 ;
      RECT 1118.5000 264.9200 1120.0000 267.9200 ;
      RECT 1114.5000 262.8250 1120.0000 264.9200 ;
      RECT 1076.5000 262.8250 1111.5000 265.8250 ;
      RECT 1060.5000 262.8250 1073.5000 265.8250 ;
      RECT 1052.3500 262.8250 1057.5000 265.8250 ;
      RECT 1044.2000 262.8250 1049.3500 265.8250 ;
      RECT 1036.0500 262.8250 1041.2000 265.8250 ;
      RECT 1027.9000 262.8250 1033.0500 265.8250 ;
      RECT 1019.7500 262.8250 1024.9000 265.8250 ;
      RECT 1011.6000 262.8250 1016.7500 265.8250 ;
      RECT 1003.4500 262.8250 1008.6000 265.8250 ;
      RECT 995.3000 262.8250 1000.4500 265.8250 ;
      RECT 987.1500 262.8250 992.3000 265.8250 ;
      RECT 979.0000 262.8250 984.1500 265.8250 ;
      RECT 970.8500 262.8250 976.0000 265.8250 ;
      RECT 962.7000 262.8250 967.8500 265.8250 ;
      RECT 954.5500 262.8250 959.7000 265.8250 ;
      RECT 946.4000 262.8250 951.5500 265.8250 ;
      RECT 938.2500 262.8250 943.4000 265.8250 ;
      RECT 930.1000 262.8250 935.2500 265.8250 ;
      RECT 921.9500 262.8250 927.1000 265.8250 ;
      RECT 913.8000 262.8250 918.9500 265.8250 ;
      RECT 905.6500 262.8250 910.8000 265.8250 ;
      RECT 897.5000 262.8250 902.6500 265.8250 ;
      RECT 889.3500 262.8250 894.5000 265.8250 ;
      RECT 881.2000 262.8250 886.3500 265.8250 ;
      RECT 873.0500 262.8250 878.2000 265.8250 ;
      RECT 864.9000 262.8250 870.0500 265.8250 ;
      RECT 856.7500 262.8250 861.9000 265.8250 ;
      RECT 848.6000 262.8250 853.7500 265.8250 ;
      RECT 840.4500 262.8250 845.6000 265.8250 ;
      RECT 832.3000 262.8250 837.4500 265.8250 ;
      RECT 824.1500 262.8250 829.3000 265.8250 ;
      RECT 816.0000 262.8250 821.1500 265.8250 ;
      RECT 807.8500 262.8250 813.0000 265.8250 ;
      RECT 799.7000 262.8250 804.8500 265.8250 ;
      RECT 791.5500 262.8250 796.7000 265.8250 ;
      RECT 783.4000 262.8250 788.5500 265.8250 ;
      RECT 775.2500 262.8250 780.4000 265.8250 ;
      RECT 767.1000 262.8250 772.2500 265.8250 ;
      RECT 758.9500 262.8250 764.1000 265.8250 ;
      RECT 750.8000 262.8250 755.9500 265.8250 ;
      RECT 742.6500 262.8250 747.8000 265.8250 ;
      RECT 734.5000 262.8250 739.6500 265.8250 ;
      RECT 726.3500 262.8250 731.5000 265.8250 ;
      RECT 718.2000 262.8250 723.3500 265.8250 ;
      RECT 710.0500 262.8250 715.2000 265.8250 ;
      RECT 701.9000 262.8250 707.0500 265.8250 ;
      RECT 693.7500 262.8250 698.9000 265.8250 ;
      RECT 685.6000 262.8250 690.7500 265.8250 ;
      RECT 677.4500 262.8250 682.6000 265.8250 ;
      RECT 669.3000 262.8250 674.4500 265.8250 ;
      RECT 661.1500 262.8250 666.3000 265.8250 ;
      RECT 653.0000 262.8250 658.1500 265.8250 ;
      RECT 644.8500 262.8250 650.0000 265.8250 ;
      RECT 636.7000 262.8250 641.8500 265.8250 ;
      RECT 628.5500 262.8250 633.7000 265.8250 ;
      RECT 620.4000 262.8250 625.5500 265.8250 ;
      RECT 612.2500 262.8250 617.4000 265.8250 ;
      RECT 604.1000 262.8250 609.2500 265.8250 ;
      RECT 595.9500 262.8250 601.1000 265.8250 ;
      RECT 587.8000 262.8250 592.9500 265.8250 ;
      RECT 579.6500 262.8250 584.8000 265.8250 ;
      RECT 571.5000 262.8250 576.6500 265.8250 ;
      RECT 563.3500 262.8250 568.5000 265.8250 ;
      RECT 555.2000 262.8250 560.3500 265.8250 ;
      RECT 547.0500 262.8250 552.2000 265.8250 ;
      RECT 538.9000 262.8250 544.0500 265.8250 ;
      RECT 530.7500 262.8250 535.9000 265.8250 ;
      RECT 522.6000 262.8250 527.7500 265.8250 ;
      RECT 514.4500 262.8250 519.6000 265.8250 ;
      RECT 506.3000 262.8250 511.4500 265.8250 ;
      RECT 498.1500 262.8250 503.3000 265.8250 ;
      RECT 490.0000 262.8250 495.1500 265.8250 ;
      RECT 481.8500 262.8250 487.0000 265.8250 ;
      RECT 473.7000 262.8250 478.8500 265.8250 ;
      RECT 465.5500 262.8250 470.7000 265.8250 ;
      RECT 457.4000 262.8250 462.5500 265.8250 ;
      RECT 449.2500 262.8250 454.4000 265.8250 ;
      RECT 441.1000 262.8250 446.2500 265.8250 ;
      RECT 432.9500 262.8250 438.1000 265.8250 ;
      RECT 424.8000 262.8250 429.9500 265.8250 ;
      RECT 416.6500 262.8250 421.8000 265.8250 ;
      RECT 396.5000 262.8250 413.6500 265.8250 ;
      RECT 346.5000 262.8250 393.5000 265.8250 ;
      RECT 326.4650 262.8250 343.5000 265.8250 ;
      RECT 317.9500 262.8250 323.4650 265.8250 ;
      RECT 309.4350 262.8250 314.9500 265.8250 ;
      RECT 300.9200 262.8250 306.4350 265.8250 ;
      RECT 292.4050 262.8250 297.9200 265.8250 ;
      RECT 283.8900 262.8250 289.4050 265.8250 ;
      RECT 275.3750 262.8250 280.8900 265.8250 ;
      RECT 266.8600 262.8250 272.3750 265.8250 ;
      RECT 258.3450 262.8250 263.8600 265.8250 ;
      RECT 249.8300 262.8250 255.3450 265.8250 ;
      RECT 241.3150 262.8250 246.8300 265.8250 ;
      RECT 232.8000 262.8250 238.3150 265.8250 ;
      RECT 224.2850 262.8250 229.8000 265.8250 ;
      RECT 215.7700 262.8250 221.2850 265.8250 ;
      RECT 207.2550 262.8250 212.7700 265.8250 ;
      RECT 198.7400 262.8250 204.2550 265.8250 ;
      RECT 190.2250 262.8250 195.7400 265.8250 ;
      RECT 181.7100 262.8250 187.2250 265.8250 ;
      RECT 173.1950 262.8250 178.7100 265.8250 ;
      RECT 164.6800 262.8250 170.1950 265.8250 ;
      RECT 156.1650 262.8250 161.6800 265.8250 ;
      RECT 147.6500 262.8250 153.1650 265.8250 ;
      RECT 139.1350 262.8250 144.6500 265.8250 ;
      RECT 130.6200 262.8250 136.1350 265.8250 ;
      RECT 122.1050 262.8250 127.6200 265.8250 ;
      RECT 113.5900 262.8250 119.1050 265.8250 ;
      RECT 105.0750 262.8250 110.5900 265.8250 ;
      RECT 96.5600 262.8250 102.0750 265.8250 ;
      RECT 88.0450 262.8250 93.5600 265.8250 ;
      RECT 79.5300 262.8250 85.0450 265.8250 ;
      RECT 71.0150 262.8250 76.5300 265.8250 ;
      RECT 62.5000 262.8250 68.0150 265.8250 ;
      RECT 46.5000 262.8250 59.5000 265.8250 ;
      RECT 8.5000 262.8250 43.5000 265.8250 ;
      RECT 0.0000 262.8250 5.5000 265.8250 ;
      RECT 0.0000 261.3000 1120.0000 262.8250 ;
      RECT 1116.6000 260.8250 1120.0000 261.3000 ;
      RECT 0.0000 258.7300 1113.6000 261.3000 ;
      RECT 1118.5000 257.8250 1120.0000 260.8250 ;
      RECT 1114.5000 255.7300 1120.0000 257.8250 ;
      RECT 1076.5000 255.7300 1111.5000 258.7300 ;
      RECT 1060.5000 255.7300 1073.5000 258.7300 ;
      RECT 1052.3500 255.7300 1057.5000 258.7300 ;
      RECT 1044.2000 255.7300 1049.3500 258.7300 ;
      RECT 1036.0500 255.7300 1041.2000 258.7300 ;
      RECT 1027.9000 255.7300 1033.0500 258.7300 ;
      RECT 1019.7500 255.7300 1024.9000 258.7300 ;
      RECT 1011.6000 255.7300 1016.7500 258.7300 ;
      RECT 1003.4500 255.7300 1008.6000 258.7300 ;
      RECT 995.3000 255.7300 1000.4500 258.7300 ;
      RECT 987.1500 255.7300 992.3000 258.7300 ;
      RECT 979.0000 255.7300 984.1500 258.7300 ;
      RECT 970.8500 255.7300 976.0000 258.7300 ;
      RECT 962.7000 255.7300 967.8500 258.7300 ;
      RECT 954.5500 255.7300 959.7000 258.7300 ;
      RECT 946.4000 255.7300 951.5500 258.7300 ;
      RECT 938.2500 255.7300 943.4000 258.7300 ;
      RECT 930.1000 255.7300 935.2500 258.7300 ;
      RECT 921.9500 255.7300 927.1000 258.7300 ;
      RECT 913.8000 255.7300 918.9500 258.7300 ;
      RECT 905.6500 255.7300 910.8000 258.7300 ;
      RECT 897.5000 255.7300 902.6500 258.7300 ;
      RECT 889.3500 255.7300 894.5000 258.7300 ;
      RECT 881.2000 255.7300 886.3500 258.7300 ;
      RECT 873.0500 255.7300 878.2000 258.7300 ;
      RECT 864.9000 255.7300 870.0500 258.7300 ;
      RECT 856.7500 255.7300 861.9000 258.7300 ;
      RECT 848.6000 255.7300 853.7500 258.7300 ;
      RECT 840.4500 255.7300 845.6000 258.7300 ;
      RECT 832.3000 255.7300 837.4500 258.7300 ;
      RECT 824.1500 255.7300 829.3000 258.7300 ;
      RECT 816.0000 255.7300 821.1500 258.7300 ;
      RECT 807.8500 255.7300 813.0000 258.7300 ;
      RECT 799.7000 255.7300 804.8500 258.7300 ;
      RECT 791.5500 255.7300 796.7000 258.7300 ;
      RECT 783.4000 255.7300 788.5500 258.7300 ;
      RECT 775.2500 255.7300 780.4000 258.7300 ;
      RECT 767.1000 255.7300 772.2500 258.7300 ;
      RECT 758.9500 255.7300 764.1000 258.7300 ;
      RECT 750.8000 255.7300 755.9500 258.7300 ;
      RECT 742.6500 255.7300 747.8000 258.7300 ;
      RECT 734.5000 255.7300 739.6500 258.7300 ;
      RECT 726.3500 255.7300 731.5000 258.7300 ;
      RECT 718.2000 255.7300 723.3500 258.7300 ;
      RECT 710.0500 255.7300 715.2000 258.7300 ;
      RECT 701.9000 255.7300 707.0500 258.7300 ;
      RECT 693.7500 255.7300 698.9000 258.7300 ;
      RECT 685.6000 255.7300 690.7500 258.7300 ;
      RECT 677.4500 255.7300 682.6000 258.7300 ;
      RECT 669.3000 255.7300 674.4500 258.7300 ;
      RECT 661.1500 255.7300 666.3000 258.7300 ;
      RECT 653.0000 255.7300 658.1500 258.7300 ;
      RECT 644.8500 255.7300 650.0000 258.7300 ;
      RECT 636.7000 255.7300 641.8500 258.7300 ;
      RECT 628.5500 255.7300 633.7000 258.7300 ;
      RECT 620.4000 255.7300 625.5500 258.7300 ;
      RECT 612.2500 255.7300 617.4000 258.7300 ;
      RECT 604.1000 255.7300 609.2500 258.7300 ;
      RECT 595.9500 255.7300 601.1000 258.7300 ;
      RECT 587.8000 255.7300 592.9500 258.7300 ;
      RECT 579.6500 255.7300 584.8000 258.7300 ;
      RECT 571.5000 255.7300 576.6500 258.7300 ;
      RECT 563.3500 255.7300 568.5000 258.7300 ;
      RECT 555.2000 255.7300 560.3500 258.7300 ;
      RECT 547.0500 255.7300 552.2000 258.7300 ;
      RECT 538.9000 255.7300 544.0500 258.7300 ;
      RECT 530.7500 255.7300 535.9000 258.7300 ;
      RECT 522.6000 255.7300 527.7500 258.7300 ;
      RECT 514.4500 255.7300 519.6000 258.7300 ;
      RECT 506.3000 255.7300 511.4500 258.7300 ;
      RECT 498.1500 255.7300 503.3000 258.7300 ;
      RECT 490.0000 255.7300 495.1500 258.7300 ;
      RECT 481.8500 255.7300 487.0000 258.7300 ;
      RECT 473.7000 255.7300 478.8500 258.7300 ;
      RECT 465.5500 255.7300 470.7000 258.7300 ;
      RECT 457.4000 255.7300 462.5500 258.7300 ;
      RECT 449.2500 255.7300 454.4000 258.7300 ;
      RECT 441.1000 255.7300 446.2500 258.7300 ;
      RECT 432.9500 255.7300 438.1000 258.7300 ;
      RECT 424.8000 255.7300 429.9500 258.7300 ;
      RECT 416.6500 255.7300 421.8000 258.7300 ;
      RECT 396.5000 255.7300 413.6500 258.7300 ;
      RECT 346.5000 255.7300 393.5000 258.7300 ;
      RECT 326.4650 255.7300 343.5000 258.7300 ;
      RECT 317.9500 255.7300 323.4650 258.7300 ;
      RECT 309.4350 255.7300 314.9500 258.7300 ;
      RECT 300.9200 255.7300 306.4350 258.7300 ;
      RECT 292.4050 255.7300 297.9200 258.7300 ;
      RECT 283.8900 255.7300 289.4050 258.7300 ;
      RECT 275.3750 255.7300 280.8900 258.7300 ;
      RECT 266.8600 255.7300 272.3750 258.7300 ;
      RECT 258.3450 255.7300 263.8600 258.7300 ;
      RECT 249.8300 255.7300 255.3450 258.7300 ;
      RECT 241.3150 255.7300 246.8300 258.7300 ;
      RECT 232.8000 255.7300 238.3150 258.7300 ;
      RECT 224.2850 255.7300 229.8000 258.7300 ;
      RECT 215.7700 255.7300 221.2850 258.7300 ;
      RECT 207.2550 255.7300 212.7700 258.7300 ;
      RECT 198.7400 255.7300 204.2550 258.7300 ;
      RECT 190.2250 255.7300 195.7400 258.7300 ;
      RECT 181.7100 255.7300 187.2250 258.7300 ;
      RECT 173.1950 255.7300 178.7100 258.7300 ;
      RECT 164.6800 255.7300 170.1950 258.7300 ;
      RECT 156.1650 255.7300 161.6800 258.7300 ;
      RECT 147.6500 255.7300 153.1650 258.7300 ;
      RECT 139.1350 255.7300 144.6500 258.7300 ;
      RECT 130.6200 255.7300 136.1350 258.7300 ;
      RECT 122.1050 255.7300 127.6200 258.7300 ;
      RECT 113.5900 255.7300 119.1050 258.7300 ;
      RECT 105.0750 255.7300 110.5900 258.7300 ;
      RECT 96.5600 255.7300 102.0750 258.7300 ;
      RECT 88.0450 255.7300 93.5600 258.7300 ;
      RECT 79.5300 255.7300 85.0450 258.7300 ;
      RECT 71.0150 255.7300 76.5300 258.7300 ;
      RECT 62.5000 255.7300 68.0150 258.7300 ;
      RECT 46.5000 255.7300 59.5000 258.7300 ;
      RECT 8.5000 255.7300 43.5000 258.7300 ;
      RECT 0.0000 255.7300 5.5000 258.7300 ;
      RECT 0.0000 254.3000 1120.0000 255.7300 ;
      RECT 1116.6000 253.7300 1120.0000 254.3000 ;
      RECT 0.0000 251.6350 1113.6000 254.3000 ;
      RECT 1118.5000 250.7300 1120.0000 253.7300 ;
      RECT 1114.5000 248.6350 1120.0000 250.7300 ;
      RECT 1076.5000 248.6350 1111.5000 251.6350 ;
      RECT 1060.5000 248.6350 1073.5000 251.6350 ;
      RECT 1052.3500 248.6350 1057.5000 251.6350 ;
      RECT 1044.2000 248.6350 1049.3500 251.6350 ;
      RECT 1036.0500 248.6350 1041.2000 251.6350 ;
      RECT 1027.9000 248.6350 1033.0500 251.6350 ;
      RECT 1019.7500 248.6350 1024.9000 251.6350 ;
      RECT 1011.6000 248.6350 1016.7500 251.6350 ;
      RECT 1003.4500 248.6350 1008.6000 251.6350 ;
      RECT 995.3000 248.6350 1000.4500 251.6350 ;
      RECT 987.1500 248.6350 992.3000 251.6350 ;
      RECT 979.0000 248.6350 984.1500 251.6350 ;
      RECT 970.8500 248.6350 976.0000 251.6350 ;
      RECT 962.7000 248.6350 967.8500 251.6350 ;
      RECT 954.5500 248.6350 959.7000 251.6350 ;
      RECT 946.4000 248.6350 951.5500 251.6350 ;
      RECT 938.2500 248.6350 943.4000 251.6350 ;
      RECT 930.1000 248.6350 935.2500 251.6350 ;
      RECT 921.9500 248.6350 927.1000 251.6350 ;
      RECT 913.8000 248.6350 918.9500 251.6350 ;
      RECT 905.6500 248.6350 910.8000 251.6350 ;
      RECT 897.5000 248.6350 902.6500 251.6350 ;
      RECT 889.3500 248.6350 894.5000 251.6350 ;
      RECT 881.2000 248.6350 886.3500 251.6350 ;
      RECT 873.0500 248.6350 878.2000 251.6350 ;
      RECT 864.9000 248.6350 870.0500 251.6350 ;
      RECT 856.7500 248.6350 861.9000 251.6350 ;
      RECT 848.6000 248.6350 853.7500 251.6350 ;
      RECT 840.4500 248.6350 845.6000 251.6350 ;
      RECT 832.3000 248.6350 837.4500 251.6350 ;
      RECT 824.1500 248.6350 829.3000 251.6350 ;
      RECT 816.0000 248.6350 821.1500 251.6350 ;
      RECT 807.8500 248.6350 813.0000 251.6350 ;
      RECT 799.7000 248.6350 804.8500 251.6350 ;
      RECT 791.5500 248.6350 796.7000 251.6350 ;
      RECT 783.4000 248.6350 788.5500 251.6350 ;
      RECT 775.2500 248.6350 780.4000 251.6350 ;
      RECT 767.1000 248.6350 772.2500 251.6350 ;
      RECT 758.9500 248.6350 764.1000 251.6350 ;
      RECT 750.8000 248.6350 755.9500 251.6350 ;
      RECT 742.6500 248.6350 747.8000 251.6350 ;
      RECT 734.5000 248.6350 739.6500 251.6350 ;
      RECT 726.3500 248.6350 731.5000 251.6350 ;
      RECT 718.2000 248.6350 723.3500 251.6350 ;
      RECT 710.0500 248.6350 715.2000 251.6350 ;
      RECT 701.9000 248.6350 707.0500 251.6350 ;
      RECT 693.7500 248.6350 698.9000 251.6350 ;
      RECT 685.6000 248.6350 690.7500 251.6350 ;
      RECT 677.4500 248.6350 682.6000 251.6350 ;
      RECT 669.3000 248.6350 674.4500 251.6350 ;
      RECT 661.1500 248.6350 666.3000 251.6350 ;
      RECT 653.0000 248.6350 658.1500 251.6350 ;
      RECT 644.8500 248.6350 650.0000 251.6350 ;
      RECT 636.7000 248.6350 641.8500 251.6350 ;
      RECT 628.5500 248.6350 633.7000 251.6350 ;
      RECT 620.4000 248.6350 625.5500 251.6350 ;
      RECT 612.2500 248.6350 617.4000 251.6350 ;
      RECT 604.1000 248.6350 609.2500 251.6350 ;
      RECT 595.9500 248.6350 601.1000 251.6350 ;
      RECT 587.8000 248.6350 592.9500 251.6350 ;
      RECT 579.6500 248.6350 584.8000 251.6350 ;
      RECT 571.5000 248.6350 576.6500 251.6350 ;
      RECT 563.3500 248.6350 568.5000 251.6350 ;
      RECT 555.2000 248.6350 560.3500 251.6350 ;
      RECT 547.0500 248.6350 552.2000 251.6350 ;
      RECT 538.9000 248.6350 544.0500 251.6350 ;
      RECT 530.7500 248.6350 535.9000 251.6350 ;
      RECT 522.6000 248.6350 527.7500 251.6350 ;
      RECT 514.4500 248.6350 519.6000 251.6350 ;
      RECT 506.3000 248.6350 511.4500 251.6350 ;
      RECT 498.1500 248.6350 503.3000 251.6350 ;
      RECT 490.0000 248.6350 495.1500 251.6350 ;
      RECT 481.8500 248.6350 487.0000 251.6350 ;
      RECT 473.7000 248.6350 478.8500 251.6350 ;
      RECT 465.5500 248.6350 470.7000 251.6350 ;
      RECT 457.4000 248.6350 462.5500 251.6350 ;
      RECT 449.2500 248.6350 454.4000 251.6350 ;
      RECT 441.1000 248.6350 446.2500 251.6350 ;
      RECT 432.9500 248.6350 438.1000 251.6350 ;
      RECT 424.8000 248.6350 429.9500 251.6350 ;
      RECT 416.6500 248.6350 421.8000 251.6350 ;
      RECT 396.5000 248.6350 413.6500 251.6350 ;
      RECT 346.5000 248.6350 393.5000 251.6350 ;
      RECT 326.4650 248.6350 343.5000 251.6350 ;
      RECT 317.9500 248.6350 323.4650 251.6350 ;
      RECT 309.4350 248.6350 314.9500 251.6350 ;
      RECT 300.9200 248.6350 306.4350 251.6350 ;
      RECT 292.4050 248.6350 297.9200 251.6350 ;
      RECT 283.8900 248.6350 289.4050 251.6350 ;
      RECT 275.3750 248.6350 280.8900 251.6350 ;
      RECT 266.8600 248.6350 272.3750 251.6350 ;
      RECT 258.3450 248.6350 263.8600 251.6350 ;
      RECT 249.8300 248.6350 255.3450 251.6350 ;
      RECT 241.3150 248.6350 246.8300 251.6350 ;
      RECT 232.8000 248.6350 238.3150 251.6350 ;
      RECT 224.2850 248.6350 229.8000 251.6350 ;
      RECT 215.7700 248.6350 221.2850 251.6350 ;
      RECT 207.2550 248.6350 212.7700 251.6350 ;
      RECT 198.7400 248.6350 204.2550 251.6350 ;
      RECT 190.2250 248.6350 195.7400 251.6350 ;
      RECT 181.7100 248.6350 187.2250 251.6350 ;
      RECT 173.1950 248.6350 178.7100 251.6350 ;
      RECT 164.6800 248.6350 170.1950 251.6350 ;
      RECT 156.1650 248.6350 161.6800 251.6350 ;
      RECT 147.6500 248.6350 153.1650 251.6350 ;
      RECT 139.1350 248.6350 144.6500 251.6350 ;
      RECT 130.6200 248.6350 136.1350 251.6350 ;
      RECT 122.1050 248.6350 127.6200 251.6350 ;
      RECT 113.5900 248.6350 119.1050 251.6350 ;
      RECT 105.0750 248.6350 110.5900 251.6350 ;
      RECT 96.5600 248.6350 102.0750 251.6350 ;
      RECT 88.0450 248.6350 93.5600 251.6350 ;
      RECT 79.5300 248.6350 85.0450 251.6350 ;
      RECT 71.0150 248.6350 76.5300 251.6350 ;
      RECT 62.5000 248.6350 68.0150 251.6350 ;
      RECT 46.5000 248.6350 59.5000 251.6350 ;
      RECT 8.5000 248.6350 43.5000 251.6350 ;
      RECT 0.0000 248.6350 5.5000 251.6350 ;
      RECT 0.0000 247.1000 1120.0000 248.6350 ;
      RECT 1116.6000 246.6350 1120.0000 247.1000 ;
      RECT 0.0000 244.5400 1113.6000 247.1000 ;
      RECT 1118.5000 243.6350 1120.0000 246.6350 ;
      RECT 1114.5000 241.5400 1120.0000 243.6350 ;
      RECT 1076.5000 241.5400 1111.5000 244.5400 ;
      RECT 1060.5000 241.5400 1073.5000 244.5400 ;
      RECT 1052.3500 241.5400 1057.5000 244.5400 ;
      RECT 1044.2000 241.5400 1049.3500 244.5400 ;
      RECT 1036.0500 241.5400 1041.2000 244.5400 ;
      RECT 1027.9000 241.5400 1033.0500 244.5400 ;
      RECT 1019.7500 241.5400 1024.9000 244.5400 ;
      RECT 1011.6000 241.5400 1016.7500 244.5400 ;
      RECT 1003.4500 241.5400 1008.6000 244.5400 ;
      RECT 995.3000 241.5400 1000.4500 244.5400 ;
      RECT 987.1500 241.5400 992.3000 244.5400 ;
      RECT 979.0000 241.5400 984.1500 244.5400 ;
      RECT 970.8500 241.5400 976.0000 244.5400 ;
      RECT 962.7000 241.5400 967.8500 244.5400 ;
      RECT 954.5500 241.5400 959.7000 244.5400 ;
      RECT 946.4000 241.5400 951.5500 244.5400 ;
      RECT 938.2500 241.5400 943.4000 244.5400 ;
      RECT 930.1000 241.5400 935.2500 244.5400 ;
      RECT 921.9500 241.5400 927.1000 244.5400 ;
      RECT 913.8000 241.5400 918.9500 244.5400 ;
      RECT 905.6500 241.5400 910.8000 244.5400 ;
      RECT 897.5000 241.5400 902.6500 244.5400 ;
      RECT 889.3500 241.5400 894.5000 244.5400 ;
      RECT 881.2000 241.5400 886.3500 244.5400 ;
      RECT 873.0500 241.5400 878.2000 244.5400 ;
      RECT 864.9000 241.5400 870.0500 244.5400 ;
      RECT 856.7500 241.5400 861.9000 244.5400 ;
      RECT 848.6000 241.5400 853.7500 244.5400 ;
      RECT 840.4500 241.5400 845.6000 244.5400 ;
      RECT 832.3000 241.5400 837.4500 244.5400 ;
      RECT 824.1500 241.5400 829.3000 244.5400 ;
      RECT 816.0000 241.5400 821.1500 244.5400 ;
      RECT 807.8500 241.5400 813.0000 244.5400 ;
      RECT 799.7000 241.5400 804.8500 244.5400 ;
      RECT 791.5500 241.5400 796.7000 244.5400 ;
      RECT 783.4000 241.5400 788.5500 244.5400 ;
      RECT 775.2500 241.5400 780.4000 244.5400 ;
      RECT 767.1000 241.5400 772.2500 244.5400 ;
      RECT 758.9500 241.5400 764.1000 244.5400 ;
      RECT 750.8000 241.5400 755.9500 244.5400 ;
      RECT 742.6500 241.5400 747.8000 244.5400 ;
      RECT 734.5000 241.5400 739.6500 244.5400 ;
      RECT 726.3500 241.5400 731.5000 244.5400 ;
      RECT 718.2000 241.5400 723.3500 244.5400 ;
      RECT 710.0500 241.5400 715.2000 244.5400 ;
      RECT 701.9000 241.5400 707.0500 244.5400 ;
      RECT 693.7500 241.5400 698.9000 244.5400 ;
      RECT 685.6000 241.5400 690.7500 244.5400 ;
      RECT 677.4500 241.5400 682.6000 244.5400 ;
      RECT 669.3000 241.5400 674.4500 244.5400 ;
      RECT 661.1500 241.5400 666.3000 244.5400 ;
      RECT 653.0000 241.5400 658.1500 244.5400 ;
      RECT 644.8500 241.5400 650.0000 244.5400 ;
      RECT 636.7000 241.5400 641.8500 244.5400 ;
      RECT 628.5500 241.5400 633.7000 244.5400 ;
      RECT 620.4000 241.5400 625.5500 244.5400 ;
      RECT 612.2500 241.5400 617.4000 244.5400 ;
      RECT 604.1000 241.5400 609.2500 244.5400 ;
      RECT 595.9500 241.5400 601.1000 244.5400 ;
      RECT 587.8000 241.5400 592.9500 244.5400 ;
      RECT 579.6500 241.5400 584.8000 244.5400 ;
      RECT 571.5000 241.5400 576.6500 244.5400 ;
      RECT 563.3500 241.5400 568.5000 244.5400 ;
      RECT 555.2000 241.5400 560.3500 244.5400 ;
      RECT 547.0500 241.5400 552.2000 244.5400 ;
      RECT 538.9000 241.5400 544.0500 244.5400 ;
      RECT 530.7500 241.5400 535.9000 244.5400 ;
      RECT 522.6000 241.5400 527.7500 244.5400 ;
      RECT 514.4500 241.5400 519.6000 244.5400 ;
      RECT 506.3000 241.5400 511.4500 244.5400 ;
      RECT 498.1500 241.5400 503.3000 244.5400 ;
      RECT 490.0000 241.5400 495.1500 244.5400 ;
      RECT 481.8500 241.5400 487.0000 244.5400 ;
      RECT 473.7000 241.5400 478.8500 244.5400 ;
      RECT 465.5500 241.5400 470.7000 244.5400 ;
      RECT 457.4000 241.5400 462.5500 244.5400 ;
      RECT 449.2500 241.5400 454.4000 244.5400 ;
      RECT 441.1000 241.5400 446.2500 244.5400 ;
      RECT 432.9500 241.5400 438.1000 244.5400 ;
      RECT 424.8000 241.5400 429.9500 244.5400 ;
      RECT 416.6500 241.5400 421.8000 244.5400 ;
      RECT 396.5000 241.5400 413.6500 244.5400 ;
      RECT 346.5000 241.5400 393.5000 244.5400 ;
      RECT 326.4650 241.5400 343.5000 244.5400 ;
      RECT 317.9500 241.5400 323.4650 244.5400 ;
      RECT 309.4350 241.5400 314.9500 244.5400 ;
      RECT 300.9200 241.5400 306.4350 244.5400 ;
      RECT 292.4050 241.5400 297.9200 244.5400 ;
      RECT 283.8900 241.5400 289.4050 244.5400 ;
      RECT 275.3750 241.5400 280.8900 244.5400 ;
      RECT 266.8600 241.5400 272.3750 244.5400 ;
      RECT 258.3450 241.5400 263.8600 244.5400 ;
      RECT 249.8300 241.5400 255.3450 244.5400 ;
      RECT 241.3150 241.5400 246.8300 244.5400 ;
      RECT 232.8000 241.5400 238.3150 244.5400 ;
      RECT 224.2850 241.5400 229.8000 244.5400 ;
      RECT 215.7700 241.5400 221.2850 244.5400 ;
      RECT 207.2550 241.5400 212.7700 244.5400 ;
      RECT 198.7400 241.5400 204.2550 244.5400 ;
      RECT 190.2250 241.5400 195.7400 244.5400 ;
      RECT 181.7100 241.5400 187.2250 244.5400 ;
      RECT 173.1950 241.5400 178.7100 244.5400 ;
      RECT 164.6800 241.5400 170.1950 244.5400 ;
      RECT 156.1650 241.5400 161.6800 244.5400 ;
      RECT 147.6500 241.5400 153.1650 244.5400 ;
      RECT 139.1350 241.5400 144.6500 244.5400 ;
      RECT 130.6200 241.5400 136.1350 244.5400 ;
      RECT 122.1050 241.5400 127.6200 244.5400 ;
      RECT 113.5900 241.5400 119.1050 244.5400 ;
      RECT 105.0750 241.5400 110.5900 244.5400 ;
      RECT 96.5600 241.5400 102.0750 244.5400 ;
      RECT 88.0450 241.5400 93.5600 244.5400 ;
      RECT 79.5300 241.5400 85.0450 244.5400 ;
      RECT 71.0150 241.5400 76.5300 244.5400 ;
      RECT 62.5000 241.5400 68.0150 244.5400 ;
      RECT 46.5000 241.5400 59.5000 244.5400 ;
      RECT 8.5000 241.5400 43.5000 244.5400 ;
      RECT 0.0000 241.5400 5.5000 244.5400 ;
      RECT 0.0000 240.1000 1120.0000 241.5400 ;
      RECT 1116.6000 239.5400 1120.0000 240.1000 ;
      RECT 0.0000 237.4450 1113.6000 240.1000 ;
      RECT 1118.5000 236.5400 1120.0000 239.5400 ;
      RECT 1114.5000 234.4450 1120.0000 236.5400 ;
      RECT 1076.5000 234.4450 1111.5000 237.4450 ;
      RECT 1060.5000 234.4450 1073.5000 237.4450 ;
      RECT 1052.3500 234.4450 1057.5000 237.4450 ;
      RECT 1044.2000 234.4450 1049.3500 237.4450 ;
      RECT 1036.0500 234.4450 1041.2000 237.4450 ;
      RECT 1027.9000 234.4450 1033.0500 237.4450 ;
      RECT 1019.7500 234.4450 1024.9000 237.4450 ;
      RECT 1011.6000 234.4450 1016.7500 237.4450 ;
      RECT 1003.4500 234.4450 1008.6000 237.4450 ;
      RECT 995.3000 234.4450 1000.4500 237.4450 ;
      RECT 987.1500 234.4450 992.3000 237.4450 ;
      RECT 979.0000 234.4450 984.1500 237.4450 ;
      RECT 970.8500 234.4450 976.0000 237.4450 ;
      RECT 962.7000 234.4450 967.8500 237.4450 ;
      RECT 954.5500 234.4450 959.7000 237.4450 ;
      RECT 946.4000 234.4450 951.5500 237.4450 ;
      RECT 938.2500 234.4450 943.4000 237.4450 ;
      RECT 930.1000 234.4450 935.2500 237.4450 ;
      RECT 921.9500 234.4450 927.1000 237.4450 ;
      RECT 913.8000 234.4450 918.9500 237.4450 ;
      RECT 905.6500 234.4450 910.8000 237.4450 ;
      RECT 897.5000 234.4450 902.6500 237.4450 ;
      RECT 889.3500 234.4450 894.5000 237.4450 ;
      RECT 881.2000 234.4450 886.3500 237.4450 ;
      RECT 873.0500 234.4450 878.2000 237.4450 ;
      RECT 864.9000 234.4450 870.0500 237.4450 ;
      RECT 856.7500 234.4450 861.9000 237.4450 ;
      RECT 848.6000 234.4450 853.7500 237.4450 ;
      RECT 840.4500 234.4450 845.6000 237.4450 ;
      RECT 832.3000 234.4450 837.4500 237.4450 ;
      RECT 824.1500 234.4450 829.3000 237.4450 ;
      RECT 816.0000 234.4450 821.1500 237.4450 ;
      RECT 807.8500 234.4450 813.0000 237.4450 ;
      RECT 799.7000 234.4450 804.8500 237.4450 ;
      RECT 791.5500 234.4450 796.7000 237.4450 ;
      RECT 783.4000 234.4450 788.5500 237.4450 ;
      RECT 775.2500 234.4450 780.4000 237.4450 ;
      RECT 767.1000 234.4450 772.2500 237.4450 ;
      RECT 758.9500 234.4450 764.1000 237.4450 ;
      RECT 750.8000 234.4450 755.9500 237.4450 ;
      RECT 742.6500 234.4450 747.8000 237.4450 ;
      RECT 734.5000 234.4450 739.6500 237.4450 ;
      RECT 726.3500 234.4450 731.5000 237.4450 ;
      RECT 718.2000 234.4450 723.3500 237.4450 ;
      RECT 710.0500 234.4450 715.2000 237.4450 ;
      RECT 701.9000 234.4450 707.0500 237.4450 ;
      RECT 693.7500 234.4450 698.9000 237.4450 ;
      RECT 685.6000 234.4450 690.7500 237.4450 ;
      RECT 677.4500 234.4450 682.6000 237.4450 ;
      RECT 669.3000 234.4450 674.4500 237.4450 ;
      RECT 661.1500 234.4450 666.3000 237.4450 ;
      RECT 653.0000 234.4450 658.1500 237.4450 ;
      RECT 644.8500 234.4450 650.0000 237.4450 ;
      RECT 636.7000 234.4450 641.8500 237.4450 ;
      RECT 628.5500 234.4450 633.7000 237.4450 ;
      RECT 620.4000 234.4450 625.5500 237.4450 ;
      RECT 612.2500 234.4450 617.4000 237.4450 ;
      RECT 604.1000 234.4450 609.2500 237.4450 ;
      RECT 595.9500 234.4450 601.1000 237.4450 ;
      RECT 587.8000 234.4450 592.9500 237.4450 ;
      RECT 579.6500 234.4450 584.8000 237.4450 ;
      RECT 571.5000 234.4450 576.6500 237.4450 ;
      RECT 563.3500 234.4450 568.5000 237.4450 ;
      RECT 555.2000 234.4450 560.3500 237.4450 ;
      RECT 547.0500 234.4450 552.2000 237.4450 ;
      RECT 538.9000 234.4450 544.0500 237.4450 ;
      RECT 530.7500 234.4450 535.9000 237.4450 ;
      RECT 522.6000 234.4450 527.7500 237.4450 ;
      RECT 514.4500 234.4450 519.6000 237.4450 ;
      RECT 506.3000 234.4450 511.4500 237.4450 ;
      RECT 498.1500 234.4450 503.3000 237.4450 ;
      RECT 490.0000 234.4450 495.1500 237.4450 ;
      RECT 481.8500 234.4450 487.0000 237.4450 ;
      RECT 473.7000 234.4450 478.8500 237.4450 ;
      RECT 465.5500 234.4450 470.7000 237.4450 ;
      RECT 457.4000 234.4450 462.5500 237.4450 ;
      RECT 449.2500 234.4450 454.4000 237.4450 ;
      RECT 441.1000 234.4450 446.2500 237.4450 ;
      RECT 432.9500 234.4450 438.1000 237.4450 ;
      RECT 424.8000 234.4450 429.9500 237.4450 ;
      RECT 416.6500 234.4450 421.8000 237.4450 ;
      RECT 396.5000 234.4450 413.6500 237.4450 ;
      RECT 346.5000 234.4450 393.5000 237.4450 ;
      RECT 326.4650 234.4450 343.5000 237.4450 ;
      RECT 317.9500 234.4450 323.4650 237.4450 ;
      RECT 309.4350 234.4450 314.9500 237.4450 ;
      RECT 300.9200 234.4450 306.4350 237.4450 ;
      RECT 292.4050 234.4450 297.9200 237.4450 ;
      RECT 283.8900 234.4450 289.4050 237.4450 ;
      RECT 275.3750 234.4450 280.8900 237.4450 ;
      RECT 266.8600 234.4450 272.3750 237.4450 ;
      RECT 258.3450 234.4450 263.8600 237.4450 ;
      RECT 249.8300 234.4450 255.3450 237.4450 ;
      RECT 241.3150 234.4450 246.8300 237.4450 ;
      RECT 232.8000 234.4450 238.3150 237.4450 ;
      RECT 224.2850 234.4450 229.8000 237.4450 ;
      RECT 215.7700 234.4450 221.2850 237.4450 ;
      RECT 207.2550 234.4450 212.7700 237.4450 ;
      RECT 198.7400 234.4450 204.2550 237.4450 ;
      RECT 190.2250 234.4450 195.7400 237.4450 ;
      RECT 181.7100 234.4450 187.2250 237.4450 ;
      RECT 173.1950 234.4450 178.7100 237.4450 ;
      RECT 164.6800 234.4450 170.1950 237.4450 ;
      RECT 156.1650 234.4450 161.6800 237.4450 ;
      RECT 147.6500 234.4450 153.1650 237.4450 ;
      RECT 139.1350 234.4450 144.6500 237.4450 ;
      RECT 130.6200 234.4450 136.1350 237.4450 ;
      RECT 122.1050 234.4450 127.6200 237.4450 ;
      RECT 113.5900 234.4450 119.1050 237.4450 ;
      RECT 105.0750 234.4450 110.5900 237.4450 ;
      RECT 96.5600 234.4450 102.0750 237.4450 ;
      RECT 88.0450 234.4450 93.5600 237.4450 ;
      RECT 79.5300 234.4450 85.0450 237.4450 ;
      RECT 71.0150 234.4450 76.5300 237.4450 ;
      RECT 62.5000 234.4450 68.0150 237.4450 ;
      RECT 46.5000 234.4450 59.5000 237.4450 ;
      RECT 8.5000 234.4450 43.5000 237.4450 ;
      RECT 0.0000 234.4450 5.5000 237.4450 ;
      RECT 0.0000 232.9000 1120.0000 234.4450 ;
      RECT 1116.6000 232.4450 1120.0000 232.9000 ;
      RECT 0.0000 230.3500 1113.6000 232.9000 ;
      RECT 1118.5000 229.4450 1120.0000 232.4450 ;
      RECT 1114.5000 227.3500 1120.0000 229.4450 ;
      RECT 1076.5000 227.3500 1111.5000 230.3500 ;
      RECT 1060.5000 227.3500 1073.5000 230.3500 ;
      RECT 1052.3500 227.3500 1057.5000 230.3500 ;
      RECT 1044.2000 227.3500 1049.3500 230.3500 ;
      RECT 1036.0500 227.3500 1041.2000 230.3500 ;
      RECT 1027.9000 227.3500 1033.0500 230.3500 ;
      RECT 1019.7500 227.3500 1024.9000 230.3500 ;
      RECT 1011.6000 227.3500 1016.7500 230.3500 ;
      RECT 1003.4500 227.3500 1008.6000 230.3500 ;
      RECT 995.3000 227.3500 1000.4500 230.3500 ;
      RECT 987.1500 227.3500 992.3000 230.3500 ;
      RECT 979.0000 227.3500 984.1500 230.3500 ;
      RECT 970.8500 227.3500 976.0000 230.3500 ;
      RECT 962.7000 227.3500 967.8500 230.3500 ;
      RECT 954.5500 227.3500 959.7000 230.3500 ;
      RECT 946.4000 227.3500 951.5500 230.3500 ;
      RECT 938.2500 227.3500 943.4000 230.3500 ;
      RECT 930.1000 227.3500 935.2500 230.3500 ;
      RECT 921.9500 227.3500 927.1000 230.3500 ;
      RECT 913.8000 227.3500 918.9500 230.3500 ;
      RECT 905.6500 227.3500 910.8000 230.3500 ;
      RECT 897.5000 227.3500 902.6500 230.3500 ;
      RECT 889.3500 227.3500 894.5000 230.3500 ;
      RECT 881.2000 227.3500 886.3500 230.3500 ;
      RECT 873.0500 227.3500 878.2000 230.3500 ;
      RECT 864.9000 227.3500 870.0500 230.3500 ;
      RECT 856.7500 227.3500 861.9000 230.3500 ;
      RECT 848.6000 227.3500 853.7500 230.3500 ;
      RECT 840.4500 227.3500 845.6000 230.3500 ;
      RECT 832.3000 227.3500 837.4500 230.3500 ;
      RECT 824.1500 227.3500 829.3000 230.3500 ;
      RECT 816.0000 227.3500 821.1500 230.3500 ;
      RECT 807.8500 227.3500 813.0000 230.3500 ;
      RECT 799.7000 227.3500 804.8500 230.3500 ;
      RECT 791.5500 227.3500 796.7000 230.3500 ;
      RECT 783.4000 227.3500 788.5500 230.3500 ;
      RECT 775.2500 227.3500 780.4000 230.3500 ;
      RECT 767.1000 227.3500 772.2500 230.3500 ;
      RECT 758.9500 227.3500 764.1000 230.3500 ;
      RECT 750.8000 227.3500 755.9500 230.3500 ;
      RECT 742.6500 227.3500 747.8000 230.3500 ;
      RECT 734.5000 227.3500 739.6500 230.3500 ;
      RECT 726.3500 227.3500 731.5000 230.3500 ;
      RECT 718.2000 227.3500 723.3500 230.3500 ;
      RECT 710.0500 227.3500 715.2000 230.3500 ;
      RECT 701.9000 227.3500 707.0500 230.3500 ;
      RECT 693.7500 227.3500 698.9000 230.3500 ;
      RECT 685.6000 227.3500 690.7500 230.3500 ;
      RECT 677.4500 227.3500 682.6000 230.3500 ;
      RECT 669.3000 227.3500 674.4500 230.3500 ;
      RECT 661.1500 227.3500 666.3000 230.3500 ;
      RECT 653.0000 227.3500 658.1500 230.3500 ;
      RECT 644.8500 227.3500 650.0000 230.3500 ;
      RECT 636.7000 227.3500 641.8500 230.3500 ;
      RECT 628.5500 227.3500 633.7000 230.3500 ;
      RECT 620.4000 227.3500 625.5500 230.3500 ;
      RECT 612.2500 227.3500 617.4000 230.3500 ;
      RECT 604.1000 227.3500 609.2500 230.3500 ;
      RECT 595.9500 227.3500 601.1000 230.3500 ;
      RECT 587.8000 227.3500 592.9500 230.3500 ;
      RECT 579.6500 227.3500 584.8000 230.3500 ;
      RECT 571.5000 227.3500 576.6500 230.3500 ;
      RECT 563.3500 227.3500 568.5000 230.3500 ;
      RECT 555.2000 227.3500 560.3500 230.3500 ;
      RECT 547.0500 227.3500 552.2000 230.3500 ;
      RECT 538.9000 227.3500 544.0500 230.3500 ;
      RECT 530.7500 227.3500 535.9000 230.3500 ;
      RECT 522.6000 227.3500 527.7500 230.3500 ;
      RECT 514.4500 227.3500 519.6000 230.3500 ;
      RECT 506.3000 227.3500 511.4500 230.3500 ;
      RECT 498.1500 227.3500 503.3000 230.3500 ;
      RECT 490.0000 227.3500 495.1500 230.3500 ;
      RECT 481.8500 227.3500 487.0000 230.3500 ;
      RECT 473.7000 227.3500 478.8500 230.3500 ;
      RECT 465.5500 227.3500 470.7000 230.3500 ;
      RECT 457.4000 227.3500 462.5500 230.3500 ;
      RECT 449.2500 227.3500 454.4000 230.3500 ;
      RECT 441.1000 227.3500 446.2500 230.3500 ;
      RECT 432.9500 227.3500 438.1000 230.3500 ;
      RECT 424.8000 227.3500 429.9500 230.3500 ;
      RECT 416.6500 227.3500 421.8000 230.3500 ;
      RECT 396.5000 227.3500 413.6500 230.3500 ;
      RECT 346.5000 227.3500 393.5000 230.3500 ;
      RECT 326.4650 227.3500 343.5000 230.3500 ;
      RECT 317.9500 227.3500 323.4650 230.3500 ;
      RECT 309.4350 227.3500 314.9500 230.3500 ;
      RECT 300.9200 227.3500 306.4350 230.3500 ;
      RECT 292.4050 227.3500 297.9200 230.3500 ;
      RECT 283.8900 227.3500 289.4050 230.3500 ;
      RECT 275.3750 227.3500 280.8900 230.3500 ;
      RECT 266.8600 227.3500 272.3750 230.3500 ;
      RECT 258.3450 227.3500 263.8600 230.3500 ;
      RECT 249.8300 227.3500 255.3450 230.3500 ;
      RECT 241.3150 227.3500 246.8300 230.3500 ;
      RECT 232.8000 227.3500 238.3150 230.3500 ;
      RECT 224.2850 227.3500 229.8000 230.3500 ;
      RECT 215.7700 227.3500 221.2850 230.3500 ;
      RECT 207.2550 227.3500 212.7700 230.3500 ;
      RECT 198.7400 227.3500 204.2550 230.3500 ;
      RECT 190.2250 227.3500 195.7400 230.3500 ;
      RECT 181.7100 227.3500 187.2250 230.3500 ;
      RECT 173.1950 227.3500 178.7100 230.3500 ;
      RECT 164.6800 227.3500 170.1950 230.3500 ;
      RECT 156.1650 227.3500 161.6800 230.3500 ;
      RECT 147.6500 227.3500 153.1650 230.3500 ;
      RECT 139.1350 227.3500 144.6500 230.3500 ;
      RECT 130.6200 227.3500 136.1350 230.3500 ;
      RECT 122.1050 227.3500 127.6200 230.3500 ;
      RECT 113.5900 227.3500 119.1050 230.3500 ;
      RECT 105.0750 227.3500 110.5900 230.3500 ;
      RECT 96.5600 227.3500 102.0750 230.3500 ;
      RECT 88.0450 227.3500 93.5600 230.3500 ;
      RECT 79.5300 227.3500 85.0450 230.3500 ;
      RECT 71.0150 227.3500 76.5300 230.3500 ;
      RECT 62.5000 227.3500 68.0150 230.3500 ;
      RECT 46.5000 227.3500 59.5000 230.3500 ;
      RECT 8.5000 227.3500 43.5000 230.3500 ;
      RECT 0.0000 227.3500 5.5000 230.3500 ;
      RECT 0.0000 225.9000 1120.0000 227.3500 ;
      RECT 1116.6000 225.3500 1120.0000 225.9000 ;
      RECT 0.0000 223.2550 1113.6000 225.9000 ;
      RECT 1118.5000 222.3500 1120.0000 225.3500 ;
      RECT 1114.5000 220.2550 1120.0000 222.3500 ;
      RECT 1076.5000 220.2550 1111.5000 223.2550 ;
      RECT 1060.5000 220.2550 1073.5000 223.2550 ;
      RECT 1052.3500 220.2550 1057.5000 223.2550 ;
      RECT 1044.2000 220.2550 1049.3500 223.2550 ;
      RECT 1036.0500 220.2550 1041.2000 223.2550 ;
      RECT 1027.9000 220.2550 1033.0500 223.2550 ;
      RECT 1019.7500 220.2550 1024.9000 223.2550 ;
      RECT 1011.6000 220.2550 1016.7500 223.2550 ;
      RECT 1003.4500 220.2550 1008.6000 223.2550 ;
      RECT 995.3000 220.2550 1000.4500 223.2550 ;
      RECT 987.1500 220.2550 992.3000 223.2550 ;
      RECT 979.0000 220.2550 984.1500 223.2550 ;
      RECT 970.8500 220.2550 976.0000 223.2550 ;
      RECT 962.7000 220.2550 967.8500 223.2550 ;
      RECT 954.5500 220.2550 959.7000 223.2550 ;
      RECT 946.4000 220.2550 951.5500 223.2550 ;
      RECT 938.2500 220.2550 943.4000 223.2550 ;
      RECT 930.1000 220.2550 935.2500 223.2550 ;
      RECT 921.9500 220.2550 927.1000 223.2550 ;
      RECT 913.8000 220.2550 918.9500 223.2550 ;
      RECT 905.6500 220.2550 910.8000 223.2550 ;
      RECT 897.5000 220.2550 902.6500 223.2550 ;
      RECT 889.3500 220.2550 894.5000 223.2550 ;
      RECT 881.2000 220.2550 886.3500 223.2550 ;
      RECT 873.0500 220.2550 878.2000 223.2550 ;
      RECT 864.9000 220.2550 870.0500 223.2550 ;
      RECT 856.7500 220.2550 861.9000 223.2550 ;
      RECT 848.6000 220.2550 853.7500 223.2550 ;
      RECT 840.4500 220.2550 845.6000 223.2550 ;
      RECT 832.3000 220.2550 837.4500 223.2550 ;
      RECT 824.1500 220.2550 829.3000 223.2550 ;
      RECT 816.0000 220.2550 821.1500 223.2550 ;
      RECT 807.8500 220.2550 813.0000 223.2550 ;
      RECT 799.7000 220.2550 804.8500 223.2550 ;
      RECT 791.5500 220.2550 796.7000 223.2550 ;
      RECT 783.4000 220.2550 788.5500 223.2550 ;
      RECT 775.2500 220.2550 780.4000 223.2550 ;
      RECT 767.1000 220.2550 772.2500 223.2550 ;
      RECT 758.9500 220.2550 764.1000 223.2550 ;
      RECT 750.8000 220.2550 755.9500 223.2550 ;
      RECT 742.6500 220.2550 747.8000 223.2550 ;
      RECT 734.5000 220.2550 739.6500 223.2550 ;
      RECT 726.3500 220.2550 731.5000 223.2550 ;
      RECT 718.2000 220.2550 723.3500 223.2550 ;
      RECT 710.0500 220.2550 715.2000 223.2550 ;
      RECT 701.9000 220.2550 707.0500 223.2550 ;
      RECT 693.7500 220.2550 698.9000 223.2550 ;
      RECT 685.6000 220.2550 690.7500 223.2550 ;
      RECT 677.4500 220.2550 682.6000 223.2550 ;
      RECT 669.3000 220.2550 674.4500 223.2550 ;
      RECT 661.1500 220.2550 666.3000 223.2550 ;
      RECT 653.0000 220.2550 658.1500 223.2550 ;
      RECT 644.8500 220.2550 650.0000 223.2550 ;
      RECT 636.7000 220.2550 641.8500 223.2550 ;
      RECT 628.5500 220.2550 633.7000 223.2550 ;
      RECT 620.4000 220.2550 625.5500 223.2550 ;
      RECT 612.2500 220.2550 617.4000 223.2550 ;
      RECT 604.1000 220.2550 609.2500 223.2550 ;
      RECT 595.9500 220.2550 601.1000 223.2550 ;
      RECT 587.8000 220.2550 592.9500 223.2550 ;
      RECT 579.6500 220.2550 584.8000 223.2550 ;
      RECT 571.5000 220.2550 576.6500 223.2550 ;
      RECT 563.3500 220.2550 568.5000 223.2550 ;
      RECT 555.2000 220.2550 560.3500 223.2550 ;
      RECT 547.0500 220.2550 552.2000 223.2550 ;
      RECT 538.9000 220.2550 544.0500 223.2550 ;
      RECT 530.7500 220.2550 535.9000 223.2550 ;
      RECT 522.6000 220.2550 527.7500 223.2550 ;
      RECT 514.4500 220.2550 519.6000 223.2550 ;
      RECT 506.3000 220.2550 511.4500 223.2550 ;
      RECT 498.1500 220.2550 503.3000 223.2550 ;
      RECT 490.0000 220.2550 495.1500 223.2550 ;
      RECT 481.8500 220.2550 487.0000 223.2550 ;
      RECT 473.7000 220.2550 478.8500 223.2550 ;
      RECT 465.5500 220.2550 470.7000 223.2550 ;
      RECT 457.4000 220.2550 462.5500 223.2550 ;
      RECT 449.2500 220.2550 454.4000 223.2550 ;
      RECT 441.1000 220.2550 446.2500 223.2550 ;
      RECT 432.9500 220.2550 438.1000 223.2550 ;
      RECT 424.8000 220.2550 429.9500 223.2550 ;
      RECT 416.6500 220.2550 421.8000 223.2550 ;
      RECT 396.5000 220.2550 413.6500 223.2550 ;
      RECT 346.5000 220.2550 393.5000 223.2550 ;
      RECT 326.4650 220.2550 343.5000 223.2550 ;
      RECT 317.9500 220.2550 323.4650 223.2550 ;
      RECT 309.4350 220.2550 314.9500 223.2550 ;
      RECT 300.9200 220.2550 306.4350 223.2550 ;
      RECT 292.4050 220.2550 297.9200 223.2550 ;
      RECT 283.8900 220.2550 289.4050 223.2550 ;
      RECT 275.3750 220.2550 280.8900 223.2550 ;
      RECT 266.8600 220.2550 272.3750 223.2550 ;
      RECT 258.3450 220.2550 263.8600 223.2550 ;
      RECT 249.8300 220.2550 255.3450 223.2550 ;
      RECT 241.3150 220.2550 246.8300 223.2550 ;
      RECT 232.8000 220.2550 238.3150 223.2550 ;
      RECT 224.2850 220.2550 229.8000 223.2550 ;
      RECT 215.7700 220.2550 221.2850 223.2550 ;
      RECT 207.2550 220.2550 212.7700 223.2550 ;
      RECT 198.7400 220.2550 204.2550 223.2550 ;
      RECT 190.2250 220.2550 195.7400 223.2550 ;
      RECT 181.7100 220.2550 187.2250 223.2550 ;
      RECT 173.1950 220.2550 178.7100 223.2550 ;
      RECT 164.6800 220.2550 170.1950 223.2550 ;
      RECT 156.1650 220.2550 161.6800 223.2550 ;
      RECT 147.6500 220.2550 153.1650 223.2550 ;
      RECT 139.1350 220.2550 144.6500 223.2550 ;
      RECT 130.6200 220.2550 136.1350 223.2550 ;
      RECT 122.1050 220.2550 127.6200 223.2550 ;
      RECT 113.5900 220.2550 119.1050 223.2550 ;
      RECT 105.0750 220.2550 110.5900 223.2550 ;
      RECT 96.5600 220.2550 102.0750 223.2550 ;
      RECT 88.0450 220.2550 93.5600 223.2550 ;
      RECT 79.5300 220.2550 85.0450 223.2550 ;
      RECT 71.0150 220.2550 76.5300 223.2550 ;
      RECT 62.5000 220.2550 68.0150 223.2550 ;
      RECT 46.5000 220.2550 59.5000 223.2550 ;
      RECT 8.5000 220.2550 43.5000 223.2550 ;
      RECT 0.0000 220.2550 5.5000 223.2550 ;
      RECT 0.0000 218.7000 1120.0000 220.2550 ;
      RECT 1116.6000 218.2550 1120.0000 218.7000 ;
      RECT 0.0000 216.1600 1113.6000 218.7000 ;
      RECT 1118.5000 215.2550 1120.0000 218.2550 ;
      RECT 1114.5000 213.1600 1120.0000 215.2550 ;
      RECT 1076.5000 213.1600 1111.5000 216.1600 ;
      RECT 1060.5000 213.1600 1073.5000 216.1600 ;
      RECT 1052.3500 213.1600 1057.5000 216.1600 ;
      RECT 1044.2000 213.1600 1049.3500 216.1600 ;
      RECT 1036.0500 213.1600 1041.2000 216.1600 ;
      RECT 1027.9000 213.1600 1033.0500 216.1600 ;
      RECT 1019.7500 213.1600 1024.9000 216.1600 ;
      RECT 1011.6000 213.1600 1016.7500 216.1600 ;
      RECT 1003.4500 213.1600 1008.6000 216.1600 ;
      RECT 995.3000 213.1600 1000.4500 216.1600 ;
      RECT 987.1500 213.1600 992.3000 216.1600 ;
      RECT 979.0000 213.1600 984.1500 216.1600 ;
      RECT 970.8500 213.1600 976.0000 216.1600 ;
      RECT 962.7000 213.1600 967.8500 216.1600 ;
      RECT 954.5500 213.1600 959.7000 216.1600 ;
      RECT 946.4000 213.1600 951.5500 216.1600 ;
      RECT 938.2500 213.1600 943.4000 216.1600 ;
      RECT 930.1000 213.1600 935.2500 216.1600 ;
      RECT 921.9500 213.1600 927.1000 216.1600 ;
      RECT 913.8000 213.1600 918.9500 216.1600 ;
      RECT 905.6500 213.1600 910.8000 216.1600 ;
      RECT 897.5000 213.1600 902.6500 216.1600 ;
      RECT 889.3500 213.1600 894.5000 216.1600 ;
      RECT 881.2000 213.1600 886.3500 216.1600 ;
      RECT 873.0500 213.1600 878.2000 216.1600 ;
      RECT 864.9000 213.1600 870.0500 216.1600 ;
      RECT 856.7500 213.1600 861.9000 216.1600 ;
      RECT 848.6000 213.1600 853.7500 216.1600 ;
      RECT 840.4500 213.1600 845.6000 216.1600 ;
      RECT 832.3000 213.1600 837.4500 216.1600 ;
      RECT 824.1500 213.1600 829.3000 216.1600 ;
      RECT 816.0000 213.1600 821.1500 216.1600 ;
      RECT 807.8500 213.1600 813.0000 216.1600 ;
      RECT 799.7000 213.1600 804.8500 216.1600 ;
      RECT 791.5500 213.1600 796.7000 216.1600 ;
      RECT 783.4000 213.1600 788.5500 216.1600 ;
      RECT 775.2500 213.1600 780.4000 216.1600 ;
      RECT 767.1000 213.1600 772.2500 216.1600 ;
      RECT 758.9500 213.1600 764.1000 216.1600 ;
      RECT 750.8000 213.1600 755.9500 216.1600 ;
      RECT 742.6500 213.1600 747.8000 216.1600 ;
      RECT 734.5000 213.1600 739.6500 216.1600 ;
      RECT 726.3500 213.1600 731.5000 216.1600 ;
      RECT 718.2000 213.1600 723.3500 216.1600 ;
      RECT 710.0500 213.1600 715.2000 216.1600 ;
      RECT 701.9000 213.1600 707.0500 216.1600 ;
      RECT 693.7500 213.1600 698.9000 216.1600 ;
      RECT 685.6000 213.1600 690.7500 216.1600 ;
      RECT 677.4500 213.1600 682.6000 216.1600 ;
      RECT 669.3000 213.1600 674.4500 216.1600 ;
      RECT 661.1500 213.1600 666.3000 216.1600 ;
      RECT 653.0000 213.1600 658.1500 216.1600 ;
      RECT 644.8500 213.1600 650.0000 216.1600 ;
      RECT 636.7000 213.1600 641.8500 216.1600 ;
      RECT 628.5500 213.1600 633.7000 216.1600 ;
      RECT 620.4000 213.1600 625.5500 216.1600 ;
      RECT 612.2500 213.1600 617.4000 216.1600 ;
      RECT 604.1000 213.1600 609.2500 216.1600 ;
      RECT 595.9500 213.1600 601.1000 216.1600 ;
      RECT 587.8000 213.1600 592.9500 216.1600 ;
      RECT 579.6500 213.1600 584.8000 216.1600 ;
      RECT 571.5000 213.1600 576.6500 216.1600 ;
      RECT 563.3500 213.1600 568.5000 216.1600 ;
      RECT 555.2000 213.1600 560.3500 216.1600 ;
      RECT 547.0500 213.1600 552.2000 216.1600 ;
      RECT 538.9000 213.1600 544.0500 216.1600 ;
      RECT 530.7500 213.1600 535.9000 216.1600 ;
      RECT 522.6000 213.1600 527.7500 216.1600 ;
      RECT 514.4500 213.1600 519.6000 216.1600 ;
      RECT 506.3000 213.1600 511.4500 216.1600 ;
      RECT 498.1500 213.1600 503.3000 216.1600 ;
      RECT 490.0000 213.1600 495.1500 216.1600 ;
      RECT 481.8500 213.1600 487.0000 216.1600 ;
      RECT 473.7000 213.1600 478.8500 216.1600 ;
      RECT 465.5500 213.1600 470.7000 216.1600 ;
      RECT 457.4000 213.1600 462.5500 216.1600 ;
      RECT 449.2500 213.1600 454.4000 216.1600 ;
      RECT 441.1000 213.1600 446.2500 216.1600 ;
      RECT 432.9500 213.1600 438.1000 216.1600 ;
      RECT 424.8000 213.1600 429.9500 216.1600 ;
      RECT 416.6500 213.1600 421.8000 216.1600 ;
      RECT 396.5000 213.1600 413.6500 216.1600 ;
      RECT 346.5000 213.1600 393.5000 216.1600 ;
      RECT 326.4650 213.1600 343.5000 216.1600 ;
      RECT 317.9500 213.1600 323.4650 216.1600 ;
      RECT 309.4350 213.1600 314.9500 216.1600 ;
      RECT 300.9200 213.1600 306.4350 216.1600 ;
      RECT 292.4050 213.1600 297.9200 216.1600 ;
      RECT 283.8900 213.1600 289.4050 216.1600 ;
      RECT 275.3750 213.1600 280.8900 216.1600 ;
      RECT 266.8600 213.1600 272.3750 216.1600 ;
      RECT 258.3450 213.1600 263.8600 216.1600 ;
      RECT 249.8300 213.1600 255.3450 216.1600 ;
      RECT 241.3150 213.1600 246.8300 216.1600 ;
      RECT 232.8000 213.1600 238.3150 216.1600 ;
      RECT 224.2850 213.1600 229.8000 216.1600 ;
      RECT 215.7700 213.1600 221.2850 216.1600 ;
      RECT 207.2550 213.1600 212.7700 216.1600 ;
      RECT 198.7400 213.1600 204.2550 216.1600 ;
      RECT 190.2250 213.1600 195.7400 216.1600 ;
      RECT 181.7100 213.1600 187.2250 216.1600 ;
      RECT 173.1950 213.1600 178.7100 216.1600 ;
      RECT 164.6800 213.1600 170.1950 216.1600 ;
      RECT 156.1650 213.1600 161.6800 216.1600 ;
      RECT 147.6500 213.1600 153.1650 216.1600 ;
      RECT 139.1350 213.1600 144.6500 216.1600 ;
      RECT 130.6200 213.1600 136.1350 216.1600 ;
      RECT 122.1050 213.1600 127.6200 216.1600 ;
      RECT 113.5900 213.1600 119.1050 216.1600 ;
      RECT 105.0750 213.1600 110.5900 216.1600 ;
      RECT 96.5600 213.1600 102.0750 216.1600 ;
      RECT 88.0450 213.1600 93.5600 216.1600 ;
      RECT 79.5300 213.1600 85.0450 216.1600 ;
      RECT 71.0150 213.1600 76.5300 216.1600 ;
      RECT 62.5000 213.1600 68.0150 216.1600 ;
      RECT 46.5000 213.1600 59.5000 216.1600 ;
      RECT 8.5000 213.1600 43.5000 216.1600 ;
      RECT 0.0000 213.1600 5.5000 216.1600 ;
      RECT 0.0000 211.7000 1120.0000 213.1600 ;
      RECT 1116.6000 211.1600 1120.0000 211.7000 ;
      RECT 0.0000 209.0650 1113.6000 211.7000 ;
      RECT 1118.5000 208.1600 1120.0000 211.1600 ;
      RECT 1114.5000 206.0650 1120.0000 208.1600 ;
      RECT 1076.5000 206.0650 1111.5000 209.0650 ;
      RECT 1060.5000 206.0650 1073.5000 209.0650 ;
      RECT 1052.3500 206.0650 1057.5000 209.0650 ;
      RECT 1044.2000 206.0650 1049.3500 209.0650 ;
      RECT 1036.0500 206.0650 1041.2000 209.0650 ;
      RECT 1027.9000 206.0650 1033.0500 209.0650 ;
      RECT 1019.7500 206.0650 1024.9000 209.0650 ;
      RECT 1011.6000 206.0650 1016.7500 209.0650 ;
      RECT 1003.4500 206.0650 1008.6000 209.0650 ;
      RECT 995.3000 206.0650 1000.4500 209.0650 ;
      RECT 987.1500 206.0650 992.3000 209.0650 ;
      RECT 979.0000 206.0650 984.1500 209.0650 ;
      RECT 970.8500 206.0650 976.0000 209.0650 ;
      RECT 962.7000 206.0650 967.8500 209.0650 ;
      RECT 954.5500 206.0650 959.7000 209.0650 ;
      RECT 946.4000 206.0650 951.5500 209.0650 ;
      RECT 938.2500 206.0650 943.4000 209.0650 ;
      RECT 930.1000 206.0650 935.2500 209.0650 ;
      RECT 921.9500 206.0650 927.1000 209.0650 ;
      RECT 913.8000 206.0650 918.9500 209.0650 ;
      RECT 905.6500 206.0650 910.8000 209.0650 ;
      RECT 897.5000 206.0650 902.6500 209.0650 ;
      RECT 889.3500 206.0650 894.5000 209.0650 ;
      RECT 881.2000 206.0650 886.3500 209.0650 ;
      RECT 873.0500 206.0650 878.2000 209.0650 ;
      RECT 864.9000 206.0650 870.0500 209.0650 ;
      RECT 856.7500 206.0650 861.9000 209.0650 ;
      RECT 848.6000 206.0650 853.7500 209.0650 ;
      RECT 840.4500 206.0650 845.6000 209.0650 ;
      RECT 832.3000 206.0650 837.4500 209.0650 ;
      RECT 824.1500 206.0650 829.3000 209.0650 ;
      RECT 816.0000 206.0650 821.1500 209.0650 ;
      RECT 807.8500 206.0650 813.0000 209.0650 ;
      RECT 799.7000 206.0650 804.8500 209.0650 ;
      RECT 791.5500 206.0650 796.7000 209.0650 ;
      RECT 783.4000 206.0650 788.5500 209.0650 ;
      RECT 775.2500 206.0650 780.4000 209.0650 ;
      RECT 767.1000 206.0650 772.2500 209.0650 ;
      RECT 758.9500 206.0650 764.1000 209.0650 ;
      RECT 750.8000 206.0650 755.9500 209.0650 ;
      RECT 742.6500 206.0650 747.8000 209.0650 ;
      RECT 734.5000 206.0650 739.6500 209.0650 ;
      RECT 726.3500 206.0650 731.5000 209.0650 ;
      RECT 718.2000 206.0650 723.3500 209.0650 ;
      RECT 710.0500 206.0650 715.2000 209.0650 ;
      RECT 701.9000 206.0650 707.0500 209.0650 ;
      RECT 693.7500 206.0650 698.9000 209.0650 ;
      RECT 685.6000 206.0650 690.7500 209.0650 ;
      RECT 677.4500 206.0650 682.6000 209.0650 ;
      RECT 669.3000 206.0650 674.4500 209.0650 ;
      RECT 661.1500 206.0650 666.3000 209.0650 ;
      RECT 653.0000 206.0650 658.1500 209.0650 ;
      RECT 644.8500 206.0650 650.0000 209.0650 ;
      RECT 636.7000 206.0650 641.8500 209.0650 ;
      RECT 628.5500 206.0650 633.7000 209.0650 ;
      RECT 620.4000 206.0650 625.5500 209.0650 ;
      RECT 612.2500 206.0650 617.4000 209.0650 ;
      RECT 604.1000 206.0650 609.2500 209.0650 ;
      RECT 595.9500 206.0650 601.1000 209.0650 ;
      RECT 587.8000 206.0650 592.9500 209.0650 ;
      RECT 579.6500 206.0650 584.8000 209.0650 ;
      RECT 571.5000 206.0650 576.6500 209.0650 ;
      RECT 563.3500 206.0650 568.5000 209.0650 ;
      RECT 555.2000 206.0650 560.3500 209.0650 ;
      RECT 547.0500 206.0650 552.2000 209.0650 ;
      RECT 538.9000 206.0650 544.0500 209.0650 ;
      RECT 530.7500 206.0650 535.9000 209.0650 ;
      RECT 522.6000 206.0650 527.7500 209.0650 ;
      RECT 514.4500 206.0650 519.6000 209.0650 ;
      RECT 506.3000 206.0650 511.4500 209.0650 ;
      RECT 498.1500 206.0650 503.3000 209.0650 ;
      RECT 490.0000 206.0650 495.1500 209.0650 ;
      RECT 481.8500 206.0650 487.0000 209.0650 ;
      RECT 473.7000 206.0650 478.8500 209.0650 ;
      RECT 465.5500 206.0650 470.7000 209.0650 ;
      RECT 457.4000 206.0650 462.5500 209.0650 ;
      RECT 449.2500 206.0650 454.4000 209.0650 ;
      RECT 441.1000 206.0650 446.2500 209.0650 ;
      RECT 432.9500 206.0650 438.1000 209.0650 ;
      RECT 424.8000 206.0650 429.9500 209.0650 ;
      RECT 416.6500 206.0650 421.8000 209.0650 ;
      RECT 396.5000 206.0650 413.6500 209.0650 ;
      RECT 346.5000 206.0650 393.5000 209.0650 ;
      RECT 326.4650 206.0650 343.5000 209.0650 ;
      RECT 317.9500 206.0650 323.4650 209.0650 ;
      RECT 309.4350 206.0650 314.9500 209.0650 ;
      RECT 300.9200 206.0650 306.4350 209.0650 ;
      RECT 292.4050 206.0650 297.9200 209.0650 ;
      RECT 283.8900 206.0650 289.4050 209.0650 ;
      RECT 275.3750 206.0650 280.8900 209.0650 ;
      RECT 266.8600 206.0650 272.3750 209.0650 ;
      RECT 258.3450 206.0650 263.8600 209.0650 ;
      RECT 249.8300 206.0650 255.3450 209.0650 ;
      RECT 241.3150 206.0650 246.8300 209.0650 ;
      RECT 232.8000 206.0650 238.3150 209.0650 ;
      RECT 224.2850 206.0650 229.8000 209.0650 ;
      RECT 215.7700 206.0650 221.2850 209.0650 ;
      RECT 207.2550 206.0650 212.7700 209.0650 ;
      RECT 198.7400 206.0650 204.2550 209.0650 ;
      RECT 190.2250 206.0650 195.7400 209.0650 ;
      RECT 181.7100 206.0650 187.2250 209.0650 ;
      RECT 173.1950 206.0650 178.7100 209.0650 ;
      RECT 164.6800 206.0650 170.1950 209.0650 ;
      RECT 156.1650 206.0650 161.6800 209.0650 ;
      RECT 147.6500 206.0650 153.1650 209.0650 ;
      RECT 139.1350 206.0650 144.6500 209.0650 ;
      RECT 130.6200 206.0650 136.1350 209.0650 ;
      RECT 122.1050 206.0650 127.6200 209.0650 ;
      RECT 113.5900 206.0650 119.1050 209.0650 ;
      RECT 105.0750 206.0650 110.5900 209.0650 ;
      RECT 96.5600 206.0650 102.0750 209.0650 ;
      RECT 88.0450 206.0650 93.5600 209.0650 ;
      RECT 79.5300 206.0650 85.0450 209.0650 ;
      RECT 71.0150 206.0650 76.5300 209.0650 ;
      RECT 62.5000 206.0650 68.0150 209.0650 ;
      RECT 46.5000 206.0650 59.5000 209.0650 ;
      RECT 8.5000 206.0650 43.5000 209.0650 ;
      RECT 0.0000 206.0650 5.5000 209.0650 ;
      RECT 0.0000 204.5000 1120.0000 206.0650 ;
      RECT 1116.6000 204.0650 1120.0000 204.5000 ;
      RECT 0.0000 201.9700 1113.6000 204.5000 ;
      RECT 1118.5000 201.0650 1120.0000 204.0650 ;
      RECT 1114.5000 198.9700 1120.0000 201.0650 ;
      RECT 1076.5000 198.9700 1111.5000 201.9700 ;
      RECT 1060.5000 198.9700 1073.5000 201.9700 ;
      RECT 1052.3500 198.9700 1057.5000 201.9700 ;
      RECT 1044.2000 198.9700 1049.3500 201.9700 ;
      RECT 1036.0500 198.9700 1041.2000 201.9700 ;
      RECT 1027.9000 198.9700 1033.0500 201.9700 ;
      RECT 1019.7500 198.9700 1024.9000 201.9700 ;
      RECT 1011.6000 198.9700 1016.7500 201.9700 ;
      RECT 1003.4500 198.9700 1008.6000 201.9700 ;
      RECT 995.3000 198.9700 1000.4500 201.9700 ;
      RECT 987.1500 198.9700 992.3000 201.9700 ;
      RECT 979.0000 198.9700 984.1500 201.9700 ;
      RECT 970.8500 198.9700 976.0000 201.9700 ;
      RECT 962.7000 198.9700 967.8500 201.9700 ;
      RECT 954.5500 198.9700 959.7000 201.9700 ;
      RECT 946.4000 198.9700 951.5500 201.9700 ;
      RECT 938.2500 198.9700 943.4000 201.9700 ;
      RECT 930.1000 198.9700 935.2500 201.9700 ;
      RECT 921.9500 198.9700 927.1000 201.9700 ;
      RECT 913.8000 198.9700 918.9500 201.9700 ;
      RECT 905.6500 198.9700 910.8000 201.9700 ;
      RECT 897.5000 198.9700 902.6500 201.9700 ;
      RECT 889.3500 198.9700 894.5000 201.9700 ;
      RECT 881.2000 198.9700 886.3500 201.9700 ;
      RECT 873.0500 198.9700 878.2000 201.9700 ;
      RECT 864.9000 198.9700 870.0500 201.9700 ;
      RECT 856.7500 198.9700 861.9000 201.9700 ;
      RECT 848.6000 198.9700 853.7500 201.9700 ;
      RECT 840.4500 198.9700 845.6000 201.9700 ;
      RECT 832.3000 198.9700 837.4500 201.9700 ;
      RECT 824.1500 198.9700 829.3000 201.9700 ;
      RECT 816.0000 198.9700 821.1500 201.9700 ;
      RECT 807.8500 198.9700 813.0000 201.9700 ;
      RECT 799.7000 198.9700 804.8500 201.9700 ;
      RECT 791.5500 198.9700 796.7000 201.9700 ;
      RECT 783.4000 198.9700 788.5500 201.9700 ;
      RECT 775.2500 198.9700 780.4000 201.9700 ;
      RECT 767.1000 198.9700 772.2500 201.9700 ;
      RECT 758.9500 198.9700 764.1000 201.9700 ;
      RECT 750.8000 198.9700 755.9500 201.9700 ;
      RECT 742.6500 198.9700 747.8000 201.9700 ;
      RECT 734.5000 198.9700 739.6500 201.9700 ;
      RECT 726.3500 198.9700 731.5000 201.9700 ;
      RECT 718.2000 198.9700 723.3500 201.9700 ;
      RECT 710.0500 198.9700 715.2000 201.9700 ;
      RECT 701.9000 198.9700 707.0500 201.9700 ;
      RECT 693.7500 198.9700 698.9000 201.9700 ;
      RECT 685.6000 198.9700 690.7500 201.9700 ;
      RECT 677.4500 198.9700 682.6000 201.9700 ;
      RECT 669.3000 198.9700 674.4500 201.9700 ;
      RECT 661.1500 198.9700 666.3000 201.9700 ;
      RECT 653.0000 198.9700 658.1500 201.9700 ;
      RECT 644.8500 198.9700 650.0000 201.9700 ;
      RECT 636.7000 198.9700 641.8500 201.9700 ;
      RECT 628.5500 198.9700 633.7000 201.9700 ;
      RECT 620.4000 198.9700 625.5500 201.9700 ;
      RECT 612.2500 198.9700 617.4000 201.9700 ;
      RECT 604.1000 198.9700 609.2500 201.9700 ;
      RECT 595.9500 198.9700 601.1000 201.9700 ;
      RECT 587.8000 198.9700 592.9500 201.9700 ;
      RECT 579.6500 198.9700 584.8000 201.9700 ;
      RECT 571.5000 198.9700 576.6500 201.9700 ;
      RECT 563.3500 198.9700 568.5000 201.9700 ;
      RECT 555.2000 198.9700 560.3500 201.9700 ;
      RECT 547.0500 198.9700 552.2000 201.9700 ;
      RECT 538.9000 198.9700 544.0500 201.9700 ;
      RECT 530.7500 198.9700 535.9000 201.9700 ;
      RECT 522.6000 198.9700 527.7500 201.9700 ;
      RECT 514.4500 198.9700 519.6000 201.9700 ;
      RECT 506.3000 198.9700 511.4500 201.9700 ;
      RECT 498.1500 198.9700 503.3000 201.9700 ;
      RECT 490.0000 198.9700 495.1500 201.9700 ;
      RECT 481.8500 198.9700 487.0000 201.9700 ;
      RECT 473.7000 198.9700 478.8500 201.9700 ;
      RECT 465.5500 198.9700 470.7000 201.9700 ;
      RECT 457.4000 198.9700 462.5500 201.9700 ;
      RECT 449.2500 198.9700 454.4000 201.9700 ;
      RECT 441.1000 198.9700 446.2500 201.9700 ;
      RECT 432.9500 198.9700 438.1000 201.9700 ;
      RECT 424.8000 198.9700 429.9500 201.9700 ;
      RECT 416.6500 198.9700 421.8000 201.9700 ;
      RECT 396.5000 198.9700 413.6500 201.9700 ;
      RECT 346.5000 198.9700 393.5000 201.9700 ;
      RECT 326.4650 198.9700 343.5000 201.9700 ;
      RECT 317.9500 198.9700 323.4650 201.9700 ;
      RECT 309.4350 198.9700 314.9500 201.9700 ;
      RECT 300.9200 198.9700 306.4350 201.9700 ;
      RECT 292.4050 198.9700 297.9200 201.9700 ;
      RECT 283.8900 198.9700 289.4050 201.9700 ;
      RECT 275.3750 198.9700 280.8900 201.9700 ;
      RECT 266.8600 198.9700 272.3750 201.9700 ;
      RECT 258.3450 198.9700 263.8600 201.9700 ;
      RECT 249.8300 198.9700 255.3450 201.9700 ;
      RECT 241.3150 198.9700 246.8300 201.9700 ;
      RECT 232.8000 198.9700 238.3150 201.9700 ;
      RECT 224.2850 198.9700 229.8000 201.9700 ;
      RECT 215.7700 198.9700 221.2850 201.9700 ;
      RECT 207.2550 198.9700 212.7700 201.9700 ;
      RECT 198.7400 198.9700 204.2550 201.9700 ;
      RECT 190.2250 198.9700 195.7400 201.9700 ;
      RECT 181.7100 198.9700 187.2250 201.9700 ;
      RECT 173.1950 198.9700 178.7100 201.9700 ;
      RECT 164.6800 198.9700 170.1950 201.9700 ;
      RECT 156.1650 198.9700 161.6800 201.9700 ;
      RECT 147.6500 198.9700 153.1650 201.9700 ;
      RECT 139.1350 198.9700 144.6500 201.9700 ;
      RECT 130.6200 198.9700 136.1350 201.9700 ;
      RECT 122.1050 198.9700 127.6200 201.9700 ;
      RECT 113.5900 198.9700 119.1050 201.9700 ;
      RECT 105.0750 198.9700 110.5900 201.9700 ;
      RECT 96.5600 198.9700 102.0750 201.9700 ;
      RECT 88.0450 198.9700 93.5600 201.9700 ;
      RECT 79.5300 198.9700 85.0450 201.9700 ;
      RECT 71.0150 198.9700 76.5300 201.9700 ;
      RECT 62.5000 198.9700 68.0150 201.9700 ;
      RECT 46.5000 198.9700 59.5000 201.9700 ;
      RECT 8.5000 198.9700 43.5000 201.9700 ;
      RECT 0.0000 198.9700 5.5000 201.9700 ;
      RECT 0.0000 197.5000 1120.0000 198.9700 ;
      RECT 1116.6000 196.9700 1120.0000 197.5000 ;
      RECT 0.0000 194.8750 1113.6000 197.5000 ;
      RECT 1118.5000 193.9700 1120.0000 196.9700 ;
      RECT 1114.5000 191.8750 1120.0000 193.9700 ;
      RECT 1076.5000 191.8750 1111.5000 194.8750 ;
      RECT 1060.5000 191.8750 1073.5000 194.8750 ;
      RECT 1052.3500 191.8750 1057.5000 194.8750 ;
      RECT 1044.2000 191.8750 1049.3500 194.8750 ;
      RECT 1036.0500 191.8750 1041.2000 194.8750 ;
      RECT 1027.9000 191.8750 1033.0500 194.8750 ;
      RECT 1019.7500 191.8750 1024.9000 194.8750 ;
      RECT 1011.6000 191.8750 1016.7500 194.8750 ;
      RECT 1003.4500 191.8750 1008.6000 194.8750 ;
      RECT 995.3000 191.8750 1000.4500 194.8750 ;
      RECT 987.1500 191.8750 992.3000 194.8750 ;
      RECT 979.0000 191.8750 984.1500 194.8750 ;
      RECT 970.8500 191.8750 976.0000 194.8750 ;
      RECT 962.7000 191.8750 967.8500 194.8750 ;
      RECT 954.5500 191.8750 959.7000 194.8750 ;
      RECT 946.4000 191.8750 951.5500 194.8750 ;
      RECT 938.2500 191.8750 943.4000 194.8750 ;
      RECT 930.1000 191.8750 935.2500 194.8750 ;
      RECT 921.9500 191.8750 927.1000 194.8750 ;
      RECT 913.8000 191.8750 918.9500 194.8750 ;
      RECT 905.6500 191.8750 910.8000 194.8750 ;
      RECT 897.5000 191.8750 902.6500 194.8750 ;
      RECT 889.3500 191.8750 894.5000 194.8750 ;
      RECT 881.2000 191.8750 886.3500 194.8750 ;
      RECT 873.0500 191.8750 878.2000 194.8750 ;
      RECT 864.9000 191.8750 870.0500 194.8750 ;
      RECT 856.7500 191.8750 861.9000 194.8750 ;
      RECT 848.6000 191.8750 853.7500 194.8750 ;
      RECT 840.4500 191.8750 845.6000 194.8750 ;
      RECT 832.3000 191.8750 837.4500 194.8750 ;
      RECT 824.1500 191.8750 829.3000 194.8750 ;
      RECT 816.0000 191.8750 821.1500 194.8750 ;
      RECT 807.8500 191.8750 813.0000 194.8750 ;
      RECT 799.7000 191.8750 804.8500 194.8750 ;
      RECT 791.5500 191.8750 796.7000 194.8750 ;
      RECT 783.4000 191.8750 788.5500 194.8750 ;
      RECT 775.2500 191.8750 780.4000 194.8750 ;
      RECT 767.1000 191.8750 772.2500 194.8750 ;
      RECT 758.9500 191.8750 764.1000 194.8750 ;
      RECT 750.8000 191.8750 755.9500 194.8750 ;
      RECT 742.6500 191.8750 747.8000 194.8750 ;
      RECT 734.5000 191.8750 739.6500 194.8750 ;
      RECT 726.3500 191.8750 731.5000 194.8750 ;
      RECT 718.2000 191.8750 723.3500 194.8750 ;
      RECT 710.0500 191.8750 715.2000 194.8750 ;
      RECT 701.9000 191.8750 707.0500 194.8750 ;
      RECT 693.7500 191.8750 698.9000 194.8750 ;
      RECT 685.6000 191.8750 690.7500 194.8750 ;
      RECT 677.4500 191.8750 682.6000 194.8750 ;
      RECT 669.3000 191.8750 674.4500 194.8750 ;
      RECT 661.1500 191.8750 666.3000 194.8750 ;
      RECT 653.0000 191.8750 658.1500 194.8750 ;
      RECT 644.8500 191.8750 650.0000 194.8750 ;
      RECT 636.7000 191.8750 641.8500 194.8750 ;
      RECT 628.5500 191.8750 633.7000 194.8750 ;
      RECT 620.4000 191.8750 625.5500 194.8750 ;
      RECT 612.2500 191.8750 617.4000 194.8750 ;
      RECT 604.1000 191.8750 609.2500 194.8750 ;
      RECT 595.9500 191.8750 601.1000 194.8750 ;
      RECT 587.8000 191.8750 592.9500 194.8750 ;
      RECT 579.6500 191.8750 584.8000 194.8750 ;
      RECT 571.5000 191.8750 576.6500 194.8750 ;
      RECT 563.3500 191.8750 568.5000 194.8750 ;
      RECT 555.2000 191.8750 560.3500 194.8750 ;
      RECT 547.0500 191.8750 552.2000 194.8750 ;
      RECT 538.9000 191.8750 544.0500 194.8750 ;
      RECT 530.7500 191.8750 535.9000 194.8750 ;
      RECT 522.6000 191.8750 527.7500 194.8750 ;
      RECT 514.4500 191.8750 519.6000 194.8750 ;
      RECT 506.3000 191.8750 511.4500 194.8750 ;
      RECT 498.1500 191.8750 503.3000 194.8750 ;
      RECT 490.0000 191.8750 495.1500 194.8750 ;
      RECT 481.8500 191.8750 487.0000 194.8750 ;
      RECT 473.7000 191.8750 478.8500 194.8750 ;
      RECT 465.5500 191.8750 470.7000 194.8750 ;
      RECT 457.4000 191.8750 462.5500 194.8750 ;
      RECT 449.2500 191.8750 454.4000 194.8750 ;
      RECT 441.1000 191.8750 446.2500 194.8750 ;
      RECT 432.9500 191.8750 438.1000 194.8750 ;
      RECT 424.8000 191.8750 429.9500 194.8750 ;
      RECT 416.6500 191.8750 421.8000 194.8750 ;
      RECT 396.5000 191.8750 413.6500 194.8750 ;
      RECT 346.5000 191.8750 393.5000 194.8750 ;
      RECT 326.4650 191.8750 343.5000 194.8750 ;
      RECT 317.9500 191.8750 323.4650 194.8750 ;
      RECT 309.4350 191.8750 314.9500 194.8750 ;
      RECT 300.9200 191.8750 306.4350 194.8750 ;
      RECT 292.4050 191.8750 297.9200 194.8750 ;
      RECT 283.8900 191.8750 289.4050 194.8750 ;
      RECT 275.3750 191.8750 280.8900 194.8750 ;
      RECT 266.8600 191.8750 272.3750 194.8750 ;
      RECT 258.3450 191.8750 263.8600 194.8750 ;
      RECT 249.8300 191.8750 255.3450 194.8750 ;
      RECT 241.3150 191.8750 246.8300 194.8750 ;
      RECT 232.8000 191.8750 238.3150 194.8750 ;
      RECT 224.2850 191.8750 229.8000 194.8750 ;
      RECT 215.7700 191.8750 221.2850 194.8750 ;
      RECT 207.2550 191.8750 212.7700 194.8750 ;
      RECT 198.7400 191.8750 204.2550 194.8750 ;
      RECT 190.2250 191.8750 195.7400 194.8750 ;
      RECT 181.7100 191.8750 187.2250 194.8750 ;
      RECT 173.1950 191.8750 178.7100 194.8750 ;
      RECT 164.6800 191.8750 170.1950 194.8750 ;
      RECT 156.1650 191.8750 161.6800 194.8750 ;
      RECT 147.6500 191.8750 153.1650 194.8750 ;
      RECT 139.1350 191.8750 144.6500 194.8750 ;
      RECT 130.6200 191.8750 136.1350 194.8750 ;
      RECT 122.1050 191.8750 127.6200 194.8750 ;
      RECT 113.5900 191.8750 119.1050 194.8750 ;
      RECT 105.0750 191.8750 110.5900 194.8750 ;
      RECT 96.5600 191.8750 102.0750 194.8750 ;
      RECT 88.0450 191.8750 93.5600 194.8750 ;
      RECT 79.5300 191.8750 85.0450 194.8750 ;
      RECT 71.0150 191.8750 76.5300 194.8750 ;
      RECT 62.5000 191.8750 68.0150 194.8750 ;
      RECT 46.5000 191.8750 59.5000 194.8750 ;
      RECT 8.5000 191.8750 43.5000 194.8750 ;
      RECT 0.0000 191.8750 5.5000 194.8750 ;
      RECT 0.0000 190.3000 1120.0000 191.8750 ;
      RECT 1116.6000 189.8750 1120.0000 190.3000 ;
      RECT 0.0000 187.7800 1113.6000 190.3000 ;
      RECT 1118.5000 186.8750 1120.0000 189.8750 ;
      RECT 1114.5000 184.7800 1120.0000 186.8750 ;
      RECT 1076.5000 184.7800 1111.5000 187.7800 ;
      RECT 1060.5000 184.7800 1073.5000 187.7800 ;
      RECT 1052.3500 184.7800 1057.5000 187.7800 ;
      RECT 1044.2000 184.7800 1049.3500 187.7800 ;
      RECT 1036.0500 184.7800 1041.2000 187.7800 ;
      RECT 1027.9000 184.7800 1033.0500 187.7800 ;
      RECT 1019.7500 184.7800 1024.9000 187.7800 ;
      RECT 1011.6000 184.7800 1016.7500 187.7800 ;
      RECT 1003.4500 184.7800 1008.6000 187.7800 ;
      RECT 995.3000 184.7800 1000.4500 187.7800 ;
      RECT 987.1500 184.7800 992.3000 187.7800 ;
      RECT 979.0000 184.7800 984.1500 187.7800 ;
      RECT 970.8500 184.7800 976.0000 187.7800 ;
      RECT 962.7000 184.7800 967.8500 187.7800 ;
      RECT 954.5500 184.7800 959.7000 187.7800 ;
      RECT 946.4000 184.7800 951.5500 187.7800 ;
      RECT 938.2500 184.7800 943.4000 187.7800 ;
      RECT 930.1000 184.7800 935.2500 187.7800 ;
      RECT 921.9500 184.7800 927.1000 187.7800 ;
      RECT 913.8000 184.7800 918.9500 187.7800 ;
      RECT 905.6500 184.7800 910.8000 187.7800 ;
      RECT 897.5000 184.7800 902.6500 187.7800 ;
      RECT 889.3500 184.7800 894.5000 187.7800 ;
      RECT 881.2000 184.7800 886.3500 187.7800 ;
      RECT 873.0500 184.7800 878.2000 187.7800 ;
      RECT 864.9000 184.7800 870.0500 187.7800 ;
      RECT 856.7500 184.7800 861.9000 187.7800 ;
      RECT 848.6000 184.7800 853.7500 187.7800 ;
      RECT 840.4500 184.7800 845.6000 187.7800 ;
      RECT 832.3000 184.7800 837.4500 187.7800 ;
      RECT 824.1500 184.7800 829.3000 187.7800 ;
      RECT 816.0000 184.7800 821.1500 187.7800 ;
      RECT 807.8500 184.7800 813.0000 187.7800 ;
      RECT 799.7000 184.7800 804.8500 187.7800 ;
      RECT 791.5500 184.7800 796.7000 187.7800 ;
      RECT 783.4000 184.7800 788.5500 187.7800 ;
      RECT 775.2500 184.7800 780.4000 187.7800 ;
      RECT 767.1000 184.7800 772.2500 187.7800 ;
      RECT 758.9500 184.7800 764.1000 187.7800 ;
      RECT 750.8000 184.7800 755.9500 187.7800 ;
      RECT 742.6500 184.7800 747.8000 187.7800 ;
      RECT 734.5000 184.7800 739.6500 187.7800 ;
      RECT 726.3500 184.7800 731.5000 187.7800 ;
      RECT 718.2000 184.7800 723.3500 187.7800 ;
      RECT 710.0500 184.7800 715.2000 187.7800 ;
      RECT 701.9000 184.7800 707.0500 187.7800 ;
      RECT 693.7500 184.7800 698.9000 187.7800 ;
      RECT 685.6000 184.7800 690.7500 187.7800 ;
      RECT 677.4500 184.7800 682.6000 187.7800 ;
      RECT 669.3000 184.7800 674.4500 187.7800 ;
      RECT 661.1500 184.7800 666.3000 187.7800 ;
      RECT 653.0000 184.7800 658.1500 187.7800 ;
      RECT 644.8500 184.7800 650.0000 187.7800 ;
      RECT 636.7000 184.7800 641.8500 187.7800 ;
      RECT 628.5500 184.7800 633.7000 187.7800 ;
      RECT 620.4000 184.7800 625.5500 187.7800 ;
      RECT 612.2500 184.7800 617.4000 187.7800 ;
      RECT 604.1000 184.7800 609.2500 187.7800 ;
      RECT 595.9500 184.7800 601.1000 187.7800 ;
      RECT 587.8000 184.7800 592.9500 187.7800 ;
      RECT 579.6500 184.7800 584.8000 187.7800 ;
      RECT 571.5000 184.7800 576.6500 187.7800 ;
      RECT 563.3500 184.7800 568.5000 187.7800 ;
      RECT 555.2000 184.7800 560.3500 187.7800 ;
      RECT 547.0500 184.7800 552.2000 187.7800 ;
      RECT 538.9000 184.7800 544.0500 187.7800 ;
      RECT 530.7500 184.7800 535.9000 187.7800 ;
      RECT 522.6000 184.7800 527.7500 187.7800 ;
      RECT 514.4500 184.7800 519.6000 187.7800 ;
      RECT 506.3000 184.7800 511.4500 187.7800 ;
      RECT 498.1500 184.7800 503.3000 187.7800 ;
      RECT 490.0000 184.7800 495.1500 187.7800 ;
      RECT 481.8500 184.7800 487.0000 187.7800 ;
      RECT 473.7000 184.7800 478.8500 187.7800 ;
      RECT 465.5500 184.7800 470.7000 187.7800 ;
      RECT 457.4000 184.7800 462.5500 187.7800 ;
      RECT 449.2500 184.7800 454.4000 187.7800 ;
      RECT 441.1000 184.7800 446.2500 187.7800 ;
      RECT 432.9500 184.7800 438.1000 187.7800 ;
      RECT 424.8000 184.7800 429.9500 187.7800 ;
      RECT 416.6500 184.7800 421.8000 187.7800 ;
      RECT 396.5000 184.7800 413.6500 187.7800 ;
      RECT 346.5000 184.7800 393.5000 187.7800 ;
      RECT 326.4650 184.7800 343.5000 187.7800 ;
      RECT 317.9500 184.7800 323.4650 187.7800 ;
      RECT 309.4350 184.7800 314.9500 187.7800 ;
      RECT 300.9200 184.7800 306.4350 187.7800 ;
      RECT 292.4050 184.7800 297.9200 187.7800 ;
      RECT 283.8900 184.7800 289.4050 187.7800 ;
      RECT 275.3750 184.7800 280.8900 187.7800 ;
      RECT 266.8600 184.7800 272.3750 187.7800 ;
      RECT 258.3450 184.7800 263.8600 187.7800 ;
      RECT 249.8300 184.7800 255.3450 187.7800 ;
      RECT 241.3150 184.7800 246.8300 187.7800 ;
      RECT 232.8000 184.7800 238.3150 187.7800 ;
      RECT 224.2850 184.7800 229.8000 187.7800 ;
      RECT 215.7700 184.7800 221.2850 187.7800 ;
      RECT 207.2550 184.7800 212.7700 187.7800 ;
      RECT 198.7400 184.7800 204.2550 187.7800 ;
      RECT 190.2250 184.7800 195.7400 187.7800 ;
      RECT 181.7100 184.7800 187.2250 187.7800 ;
      RECT 173.1950 184.7800 178.7100 187.7800 ;
      RECT 164.6800 184.7800 170.1950 187.7800 ;
      RECT 156.1650 184.7800 161.6800 187.7800 ;
      RECT 147.6500 184.7800 153.1650 187.7800 ;
      RECT 139.1350 184.7800 144.6500 187.7800 ;
      RECT 130.6200 184.7800 136.1350 187.7800 ;
      RECT 122.1050 184.7800 127.6200 187.7800 ;
      RECT 113.5900 184.7800 119.1050 187.7800 ;
      RECT 105.0750 184.7800 110.5900 187.7800 ;
      RECT 96.5600 184.7800 102.0750 187.7800 ;
      RECT 88.0450 184.7800 93.5600 187.7800 ;
      RECT 79.5300 184.7800 85.0450 187.7800 ;
      RECT 71.0150 184.7800 76.5300 187.7800 ;
      RECT 62.5000 184.7800 68.0150 187.7800 ;
      RECT 46.5000 184.7800 59.5000 187.7800 ;
      RECT 8.5000 184.7800 43.5000 187.7800 ;
      RECT 0.0000 184.7800 5.5000 187.7800 ;
      RECT 0.0000 183.3000 1120.0000 184.7800 ;
      RECT 1116.6000 182.7800 1120.0000 183.3000 ;
      RECT 0.0000 180.6850 1113.6000 183.3000 ;
      RECT 1118.5000 179.7800 1120.0000 182.7800 ;
      RECT 1114.5000 177.6850 1120.0000 179.7800 ;
      RECT 1076.5000 177.6850 1111.5000 180.6850 ;
      RECT 1060.5000 177.6850 1073.5000 180.6850 ;
      RECT 1052.3500 177.6850 1057.5000 180.6850 ;
      RECT 1044.2000 177.6850 1049.3500 180.6850 ;
      RECT 1036.0500 177.6850 1041.2000 180.6850 ;
      RECT 1027.9000 177.6850 1033.0500 180.6850 ;
      RECT 1019.7500 177.6850 1024.9000 180.6850 ;
      RECT 1011.6000 177.6850 1016.7500 180.6850 ;
      RECT 1003.4500 177.6850 1008.6000 180.6850 ;
      RECT 995.3000 177.6850 1000.4500 180.6850 ;
      RECT 987.1500 177.6850 992.3000 180.6850 ;
      RECT 979.0000 177.6850 984.1500 180.6850 ;
      RECT 970.8500 177.6850 976.0000 180.6850 ;
      RECT 962.7000 177.6850 967.8500 180.6850 ;
      RECT 954.5500 177.6850 959.7000 180.6850 ;
      RECT 946.4000 177.6850 951.5500 180.6850 ;
      RECT 938.2500 177.6850 943.4000 180.6850 ;
      RECT 930.1000 177.6850 935.2500 180.6850 ;
      RECT 921.9500 177.6850 927.1000 180.6850 ;
      RECT 913.8000 177.6850 918.9500 180.6850 ;
      RECT 905.6500 177.6850 910.8000 180.6850 ;
      RECT 897.5000 177.6850 902.6500 180.6850 ;
      RECT 889.3500 177.6850 894.5000 180.6850 ;
      RECT 881.2000 177.6850 886.3500 180.6850 ;
      RECT 873.0500 177.6850 878.2000 180.6850 ;
      RECT 864.9000 177.6850 870.0500 180.6850 ;
      RECT 856.7500 177.6850 861.9000 180.6850 ;
      RECT 848.6000 177.6850 853.7500 180.6850 ;
      RECT 840.4500 177.6850 845.6000 180.6850 ;
      RECT 832.3000 177.6850 837.4500 180.6850 ;
      RECT 824.1500 177.6850 829.3000 180.6850 ;
      RECT 816.0000 177.6850 821.1500 180.6850 ;
      RECT 807.8500 177.6850 813.0000 180.6850 ;
      RECT 799.7000 177.6850 804.8500 180.6850 ;
      RECT 791.5500 177.6850 796.7000 180.6850 ;
      RECT 783.4000 177.6850 788.5500 180.6850 ;
      RECT 775.2500 177.6850 780.4000 180.6850 ;
      RECT 767.1000 177.6850 772.2500 180.6850 ;
      RECT 758.9500 177.6850 764.1000 180.6850 ;
      RECT 750.8000 177.6850 755.9500 180.6850 ;
      RECT 742.6500 177.6850 747.8000 180.6850 ;
      RECT 734.5000 177.6850 739.6500 180.6850 ;
      RECT 726.3500 177.6850 731.5000 180.6850 ;
      RECT 718.2000 177.6850 723.3500 180.6850 ;
      RECT 710.0500 177.6850 715.2000 180.6850 ;
      RECT 701.9000 177.6850 707.0500 180.6850 ;
      RECT 693.7500 177.6850 698.9000 180.6850 ;
      RECT 685.6000 177.6850 690.7500 180.6850 ;
      RECT 677.4500 177.6850 682.6000 180.6850 ;
      RECT 669.3000 177.6850 674.4500 180.6850 ;
      RECT 661.1500 177.6850 666.3000 180.6850 ;
      RECT 653.0000 177.6850 658.1500 180.6850 ;
      RECT 644.8500 177.6850 650.0000 180.6850 ;
      RECT 636.7000 177.6850 641.8500 180.6850 ;
      RECT 628.5500 177.6850 633.7000 180.6850 ;
      RECT 620.4000 177.6850 625.5500 180.6850 ;
      RECT 612.2500 177.6850 617.4000 180.6850 ;
      RECT 604.1000 177.6850 609.2500 180.6850 ;
      RECT 595.9500 177.6850 601.1000 180.6850 ;
      RECT 587.8000 177.6850 592.9500 180.6850 ;
      RECT 579.6500 177.6850 584.8000 180.6850 ;
      RECT 571.5000 177.6850 576.6500 180.6850 ;
      RECT 563.3500 177.6850 568.5000 180.6850 ;
      RECT 555.2000 177.6850 560.3500 180.6850 ;
      RECT 547.0500 177.6850 552.2000 180.6850 ;
      RECT 538.9000 177.6850 544.0500 180.6850 ;
      RECT 530.7500 177.6850 535.9000 180.6850 ;
      RECT 522.6000 177.6850 527.7500 180.6850 ;
      RECT 514.4500 177.6850 519.6000 180.6850 ;
      RECT 506.3000 177.6850 511.4500 180.6850 ;
      RECT 498.1500 177.6850 503.3000 180.6850 ;
      RECT 490.0000 177.6850 495.1500 180.6850 ;
      RECT 481.8500 177.6850 487.0000 180.6850 ;
      RECT 473.7000 177.6850 478.8500 180.6850 ;
      RECT 465.5500 177.6850 470.7000 180.6850 ;
      RECT 457.4000 177.6850 462.5500 180.6850 ;
      RECT 449.2500 177.6850 454.4000 180.6850 ;
      RECT 441.1000 177.6850 446.2500 180.6850 ;
      RECT 432.9500 177.6850 438.1000 180.6850 ;
      RECT 424.8000 177.6850 429.9500 180.6850 ;
      RECT 416.6500 177.6850 421.8000 180.6850 ;
      RECT 396.5000 177.6850 413.6500 180.6850 ;
      RECT 346.5000 177.6850 393.5000 180.6850 ;
      RECT 326.4650 177.6850 343.5000 180.6850 ;
      RECT 317.9500 177.6850 323.4650 180.6850 ;
      RECT 309.4350 177.6850 314.9500 180.6850 ;
      RECT 300.9200 177.6850 306.4350 180.6850 ;
      RECT 292.4050 177.6850 297.9200 180.6850 ;
      RECT 283.8900 177.6850 289.4050 180.6850 ;
      RECT 275.3750 177.6850 280.8900 180.6850 ;
      RECT 266.8600 177.6850 272.3750 180.6850 ;
      RECT 258.3450 177.6850 263.8600 180.6850 ;
      RECT 249.8300 177.6850 255.3450 180.6850 ;
      RECT 241.3150 177.6850 246.8300 180.6850 ;
      RECT 232.8000 177.6850 238.3150 180.6850 ;
      RECT 224.2850 177.6850 229.8000 180.6850 ;
      RECT 215.7700 177.6850 221.2850 180.6850 ;
      RECT 207.2550 177.6850 212.7700 180.6850 ;
      RECT 198.7400 177.6850 204.2550 180.6850 ;
      RECT 190.2250 177.6850 195.7400 180.6850 ;
      RECT 181.7100 177.6850 187.2250 180.6850 ;
      RECT 173.1950 177.6850 178.7100 180.6850 ;
      RECT 164.6800 177.6850 170.1950 180.6850 ;
      RECT 156.1650 177.6850 161.6800 180.6850 ;
      RECT 147.6500 177.6850 153.1650 180.6850 ;
      RECT 139.1350 177.6850 144.6500 180.6850 ;
      RECT 130.6200 177.6850 136.1350 180.6850 ;
      RECT 122.1050 177.6850 127.6200 180.6850 ;
      RECT 113.5900 177.6850 119.1050 180.6850 ;
      RECT 105.0750 177.6850 110.5900 180.6850 ;
      RECT 96.5600 177.6850 102.0750 180.6850 ;
      RECT 88.0450 177.6850 93.5600 180.6850 ;
      RECT 79.5300 177.6850 85.0450 180.6850 ;
      RECT 71.0150 177.6850 76.5300 180.6850 ;
      RECT 62.5000 177.6850 68.0150 180.6850 ;
      RECT 46.5000 177.6850 59.5000 180.6850 ;
      RECT 8.5000 177.6850 43.5000 180.6850 ;
      RECT 0.0000 177.6850 5.5000 180.6850 ;
      RECT 0.0000 176.1000 1120.0000 177.6850 ;
      RECT 1116.6000 175.6850 1120.0000 176.1000 ;
      RECT 0.0000 173.5900 1113.6000 176.1000 ;
      RECT 1118.5000 172.6850 1120.0000 175.6850 ;
      RECT 1114.5000 170.5900 1120.0000 172.6850 ;
      RECT 1076.5000 170.5900 1111.5000 173.5900 ;
      RECT 1060.5000 170.5900 1073.5000 173.5900 ;
      RECT 1052.3500 170.5900 1057.5000 173.5900 ;
      RECT 1044.2000 170.5900 1049.3500 173.5900 ;
      RECT 1036.0500 170.5900 1041.2000 173.5900 ;
      RECT 1027.9000 170.5900 1033.0500 173.5900 ;
      RECT 1019.7500 170.5900 1024.9000 173.5900 ;
      RECT 1011.6000 170.5900 1016.7500 173.5900 ;
      RECT 1003.4500 170.5900 1008.6000 173.5900 ;
      RECT 995.3000 170.5900 1000.4500 173.5900 ;
      RECT 987.1500 170.5900 992.3000 173.5900 ;
      RECT 979.0000 170.5900 984.1500 173.5900 ;
      RECT 970.8500 170.5900 976.0000 173.5900 ;
      RECT 962.7000 170.5900 967.8500 173.5900 ;
      RECT 954.5500 170.5900 959.7000 173.5900 ;
      RECT 946.4000 170.5900 951.5500 173.5900 ;
      RECT 938.2500 170.5900 943.4000 173.5900 ;
      RECT 930.1000 170.5900 935.2500 173.5900 ;
      RECT 921.9500 170.5900 927.1000 173.5900 ;
      RECT 913.8000 170.5900 918.9500 173.5900 ;
      RECT 905.6500 170.5900 910.8000 173.5900 ;
      RECT 897.5000 170.5900 902.6500 173.5900 ;
      RECT 889.3500 170.5900 894.5000 173.5900 ;
      RECT 881.2000 170.5900 886.3500 173.5900 ;
      RECT 873.0500 170.5900 878.2000 173.5900 ;
      RECT 864.9000 170.5900 870.0500 173.5900 ;
      RECT 856.7500 170.5900 861.9000 173.5900 ;
      RECT 848.6000 170.5900 853.7500 173.5900 ;
      RECT 840.4500 170.5900 845.6000 173.5900 ;
      RECT 832.3000 170.5900 837.4500 173.5900 ;
      RECT 824.1500 170.5900 829.3000 173.5900 ;
      RECT 816.0000 170.5900 821.1500 173.5900 ;
      RECT 807.8500 170.5900 813.0000 173.5900 ;
      RECT 799.7000 170.5900 804.8500 173.5900 ;
      RECT 791.5500 170.5900 796.7000 173.5900 ;
      RECT 783.4000 170.5900 788.5500 173.5900 ;
      RECT 775.2500 170.5900 780.4000 173.5900 ;
      RECT 767.1000 170.5900 772.2500 173.5900 ;
      RECT 758.9500 170.5900 764.1000 173.5900 ;
      RECT 750.8000 170.5900 755.9500 173.5900 ;
      RECT 742.6500 170.5900 747.8000 173.5900 ;
      RECT 734.5000 170.5900 739.6500 173.5900 ;
      RECT 726.3500 170.5900 731.5000 173.5900 ;
      RECT 718.2000 170.5900 723.3500 173.5900 ;
      RECT 710.0500 170.5900 715.2000 173.5900 ;
      RECT 701.9000 170.5900 707.0500 173.5900 ;
      RECT 693.7500 170.5900 698.9000 173.5900 ;
      RECT 685.6000 170.5900 690.7500 173.5900 ;
      RECT 677.4500 170.5900 682.6000 173.5900 ;
      RECT 669.3000 170.5900 674.4500 173.5900 ;
      RECT 661.1500 170.5900 666.3000 173.5900 ;
      RECT 653.0000 170.5900 658.1500 173.5900 ;
      RECT 644.8500 170.5900 650.0000 173.5900 ;
      RECT 636.7000 170.5900 641.8500 173.5900 ;
      RECT 628.5500 170.5900 633.7000 173.5900 ;
      RECT 620.4000 170.5900 625.5500 173.5900 ;
      RECT 612.2500 170.5900 617.4000 173.5900 ;
      RECT 604.1000 170.5900 609.2500 173.5900 ;
      RECT 595.9500 170.5900 601.1000 173.5900 ;
      RECT 587.8000 170.5900 592.9500 173.5900 ;
      RECT 579.6500 170.5900 584.8000 173.5900 ;
      RECT 571.5000 170.5900 576.6500 173.5900 ;
      RECT 563.3500 170.5900 568.5000 173.5900 ;
      RECT 555.2000 170.5900 560.3500 173.5900 ;
      RECT 547.0500 170.5900 552.2000 173.5900 ;
      RECT 538.9000 170.5900 544.0500 173.5900 ;
      RECT 530.7500 170.5900 535.9000 173.5900 ;
      RECT 522.6000 170.5900 527.7500 173.5900 ;
      RECT 514.4500 170.5900 519.6000 173.5900 ;
      RECT 506.3000 170.5900 511.4500 173.5900 ;
      RECT 498.1500 170.5900 503.3000 173.5900 ;
      RECT 490.0000 170.5900 495.1500 173.5900 ;
      RECT 481.8500 170.5900 487.0000 173.5900 ;
      RECT 473.7000 170.5900 478.8500 173.5900 ;
      RECT 465.5500 170.5900 470.7000 173.5900 ;
      RECT 457.4000 170.5900 462.5500 173.5900 ;
      RECT 449.2500 170.5900 454.4000 173.5900 ;
      RECT 441.1000 170.5900 446.2500 173.5900 ;
      RECT 432.9500 170.5900 438.1000 173.5900 ;
      RECT 424.8000 170.5900 429.9500 173.5900 ;
      RECT 416.6500 170.5900 421.8000 173.5900 ;
      RECT 396.5000 170.5900 413.6500 173.5900 ;
      RECT 346.5000 170.5900 393.5000 173.5900 ;
      RECT 326.4650 170.5900 343.5000 173.5900 ;
      RECT 317.9500 170.5900 323.4650 173.5900 ;
      RECT 309.4350 170.5900 314.9500 173.5900 ;
      RECT 300.9200 170.5900 306.4350 173.5900 ;
      RECT 292.4050 170.5900 297.9200 173.5900 ;
      RECT 283.8900 170.5900 289.4050 173.5900 ;
      RECT 275.3750 170.5900 280.8900 173.5900 ;
      RECT 266.8600 170.5900 272.3750 173.5900 ;
      RECT 258.3450 170.5900 263.8600 173.5900 ;
      RECT 249.8300 170.5900 255.3450 173.5900 ;
      RECT 241.3150 170.5900 246.8300 173.5900 ;
      RECT 232.8000 170.5900 238.3150 173.5900 ;
      RECT 224.2850 170.5900 229.8000 173.5900 ;
      RECT 215.7700 170.5900 221.2850 173.5900 ;
      RECT 207.2550 170.5900 212.7700 173.5900 ;
      RECT 198.7400 170.5900 204.2550 173.5900 ;
      RECT 190.2250 170.5900 195.7400 173.5900 ;
      RECT 181.7100 170.5900 187.2250 173.5900 ;
      RECT 173.1950 170.5900 178.7100 173.5900 ;
      RECT 164.6800 170.5900 170.1950 173.5900 ;
      RECT 156.1650 170.5900 161.6800 173.5900 ;
      RECT 147.6500 170.5900 153.1650 173.5900 ;
      RECT 139.1350 170.5900 144.6500 173.5900 ;
      RECT 130.6200 170.5900 136.1350 173.5900 ;
      RECT 122.1050 170.5900 127.6200 173.5900 ;
      RECT 113.5900 170.5900 119.1050 173.5900 ;
      RECT 105.0750 170.5900 110.5900 173.5900 ;
      RECT 96.5600 170.5900 102.0750 173.5900 ;
      RECT 88.0450 170.5900 93.5600 173.5900 ;
      RECT 79.5300 170.5900 85.0450 173.5900 ;
      RECT 71.0150 170.5900 76.5300 173.5900 ;
      RECT 62.5000 170.5900 68.0150 173.5900 ;
      RECT 46.5000 170.5900 59.5000 173.5900 ;
      RECT 8.5000 170.5900 43.5000 173.5900 ;
      RECT 0.0000 170.5900 5.5000 173.5900 ;
      RECT 0.0000 169.1000 1120.0000 170.5900 ;
      RECT 1116.6000 168.5900 1120.0000 169.1000 ;
      RECT 0.0000 166.4950 1113.6000 169.1000 ;
      RECT 1118.5000 165.5900 1120.0000 168.5900 ;
      RECT 1114.5000 163.4950 1120.0000 165.5900 ;
      RECT 1076.5000 163.4950 1111.5000 166.4950 ;
      RECT 1060.5000 163.4950 1073.5000 166.4950 ;
      RECT 1052.3500 163.4950 1057.5000 166.4950 ;
      RECT 1044.2000 163.4950 1049.3500 166.4950 ;
      RECT 1036.0500 163.4950 1041.2000 166.4950 ;
      RECT 1027.9000 163.4950 1033.0500 166.4950 ;
      RECT 1019.7500 163.4950 1024.9000 166.4950 ;
      RECT 1011.6000 163.4950 1016.7500 166.4950 ;
      RECT 1003.4500 163.4950 1008.6000 166.4950 ;
      RECT 995.3000 163.4950 1000.4500 166.4950 ;
      RECT 987.1500 163.4950 992.3000 166.4950 ;
      RECT 979.0000 163.4950 984.1500 166.4950 ;
      RECT 970.8500 163.4950 976.0000 166.4950 ;
      RECT 962.7000 163.4950 967.8500 166.4950 ;
      RECT 954.5500 163.4950 959.7000 166.4950 ;
      RECT 946.4000 163.4950 951.5500 166.4950 ;
      RECT 938.2500 163.4950 943.4000 166.4950 ;
      RECT 930.1000 163.4950 935.2500 166.4950 ;
      RECT 921.9500 163.4950 927.1000 166.4950 ;
      RECT 913.8000 163.4950 918.9500 166.4950 ;
      RECT 905.6500 163.4950 910.8000 166.4950 ;
      RECT 897.5000 163.4950 902.6500 166.4950 ;
      RECT 889.3500 163.4950 894.5000 166.4950 ;
      RECT 881.2000 163.4950 886.3500 166.4950 ;
      RECT 873.0500 163.4950 878.2000 166.4950 ;
      RECT 864.9000 163.4950 870.0500 166.4950 ;
      RECT 856.7500 163.4950 861.9000 166.4950 ;
      RECT 848.6000 163.4950 853.7500 166.4950 ;
      RECT 840.4500 163.4950 845.6000 166.4950 ;
      RECT 832.3000 163.4950 837.4500 166.4950 ;
      RECT 824.1500 163.4950 829.3000 166.4950 ;
      RECT 816.0000 163.4950 821.1500 166.4950 ;
      RECT 807.8500 163.4950 813.0000 166.4950 ;
      RECT 799.7000 163.4950 804.8500 166.4950 ;
      RECT 791.5500 163.4950 796.7000 166.4950 ;
      RECT 783.4000 163.4950 788.5500 166.4950 ;
      RECT 775.2500 163.4950 780.4000 166.4950 ;
      RECT 767.1000 163.4950 772.2500 166.4950 ;
      RECT 758.9500 163.4950 764.1000 166.4950 ;
      RECT 750.8000 163.4950 755.9500 166.4950 ;
      RECT 742.6500 163.4950 747.8000 166.4950 ;
      RECT 734.5000 163.4950 739.6500 166.4950 ;
      RECT 726.3500 163.4950 731.5000 166.4950 ;
      RECT 718.2000 163.4950 723.3500 166.4950 ;
      RECT 710.0500 163.4950 715.2000 166.4950 ;
      RECT 701.9000 163.4950 707.0500 166.4950 ;
      RECT 693.7500 163.4950 698.9000 166.4950 ;
      RECT 685.6000 163.4950 690.7500 166.4950 ;
      RECT 677.4500 163.4950 682.6000 166.4950 ;
      RECT 669.3000 163.4950 674.4500 166.4950 ;
      RECT 661.1500 163.4950 666.3000 166.4950 ;
      RECT 653.0000 163.4950 658.1500 166.4950 ;
      RECT 644.8500 163.4950 650.0000 166.4950 ;
      RECT 636.7000 163.4950 641.8500 166.4950 ;
      RECT 628.5500 163.4950 633.7000 166.4950 ;
      RECT 620.4000 163.4950 625.5500 166.4950 ;
      RECT 612.2500 163.4950 617.4000 166.4950 ;
      RECT 604.1000 163.4950 609.2500 166.4950 ;
      RECT 595.9500 163.4950 601.1000 166.4950 ;
      RECT 587.8000 163.4950 592.9500 166.4950 ;
      RECT 579.6500 163.4950 584.8000 166.4950 ;
      RECT 571.5000 163.4950 576.6500 166.4950 ;
      RECT 563.3500 163.4950 568.5000 166.4950 ;
      RECT 555.2000 163.4950 560.3500 166.4950 ;
      RECT 547.0500 163.4950 552.2000 166.4950 ;
      RECT 538.9000 163.4950 544.0500 166.4950 ;
      RECT 530.7500 163.4950 535.9000 166.4950 ;
      RECT 522.6000 163.4950 527.7500 166.4950 ;
      RECT 514.4500 163.4950 519.6000 166.4950 ;
      RECT 506.3000 163.4950 511.4500 166.4950 ;
      RECT 498.1500 163.4950 503.3000 166.4950 ;
      RECT 490.0000 163.4950 495.1500 166.4950 ;
      RECT 481.8500 163.4950 487.0000 166.4950 ;
      RECT 473.7000 163.4950 478.8500 166.4950 ;
      RECT 465.5500 163.4950 470.7000 166.4950 ;
      RECT 457.4000 163.4950 462.5500 166.4950 ;
      RECT 449.2500 163.4950 454.4000 166.4950 ;
      RECT 441.1000 163.4950 446.2500 166.4950 ;
      RECT 432.9500 163.4950 438.1000 166.4950 ;
      RECT 424.8000 163.4950 429.9500 166.4950 ;
      RECT 416.6500 163.4950 421.8000 166.4950 ;
      RECT 396.5000 163.4950 413.6500 166.4950 ;
      RECT 346.5000 163.4950 393.5000 166.4950 ;
      RECT 326.4650 163.4950 343.5000 166.4950 ;
      RECT 317.9500 163.4950 323.4650 166.4950 ;
      RECT 309.4350 163.4950 314.9500 166.4950 ;
      RECT 300.9200 163.4950 306.4350 166.4950 ;
      RECT 292.4050 163.4950 297.9200 166.4950 ;
      RECT 283.8900 163.4950 289.4050 166.4950 ;
      RECT 275.3750 163.4950 280.8900 166.4950 ;
      RECT 266.8600 163.4950 272.3750 166.4950 ;
      RECT 258.3450 163.4950 263.8600 166.4950 ;
      RECT 249.8300 163.4950 255.3450 166.4950 ;
      RECT 241.3150 163.4950 246.8300 166.4950 ;
      RECT 232.8000 163.4950 238.3150 166.4950 ;
      RECT 224.2850 163.4950 229.8000 166.4950 ;
      RECT 215.7700 163.4950 221.2850 166.4950 ;
      RECT 207.2550 163.4950 212.7700 166.4950 ;
      RECT 198.7400 163.4950 204.2550 166.4950 ;
      RECT 190.2250 163.4950 195.7400 166.4950 ;
      RECT 181.7100 163.4950 187.2250 166.4950 ;
      RECT 173.1950 163.4950 178.7100 166.4950 ;
      RECT 164.6800 163.4950 170.1950 166.4950 ;
      RECT 156.1650 163.4950 161.6800 166.4950 ;
      RECT 147.6500 163.4950 153.1650 166.4950 ;
      RECT 139.1350 163.4950 144.6500 166.4950 ;
      RECT 130.6200 163.4950 136.1350 166.4950 ;
      RECT 122.1050 163.4950 127.6200 166.4950 ;
      RECT 113.5900 163.4950 119.1050 166.4950 ;
      RECT 105.0750 163.4950 110.5900 166.4950 ;
      RECT 96.5600 163.4950 102.0750 166.4950 ;
      RECT 88.0450 163.4950 93.5600 166.4950 ;
      RECT 79.5300 163.4950 85.0450 166.4950 ;
      RECT 71.0150 163.4950 76.5300 166.4950 ;
      RECT 62.5000 163.4950 68.0150 166.4950 ;
      RECT 46.5000 163.4950 59.5000 166.4950 ;
      RECT 8.5000 163.4950 43.5000 166.4950 ;
      RECT 0.0000 163.4950 5.5000 166.4950 ;
      RECT 0.0000 161.9000 1120.0000 163.4950 ;
      RECT 1116.6000 161.4950 1120.0000 161.9000 ;
      RECT 0.0000 159.4000 1113.6000 161.9000 ;
      RECT 1118.5000 158.4950 1120.0000 161.4950 ;
      RECT 1114.5000 156.4000 1120.0000 158.4950 ;
      RECT 1076.5000 156.4000 1111.5000 159.4000 ;
      RECT 1060.5000 156.4000 1073.5000 159.4000 ;
      RECT 1052.3500 156.4000 1057.5000 159.4000 ;
      RECT 1044.2000 156.4000 1049.3500 159.4000 ;
      RECT 1036.0500 156.4000 1041.2000 159.4000 ;
      RECT 1027.9000 156.4000 1033.0500 159.4000 ;
      RECT 1019.7500 156.4000 1024.9000 159.4000 ;
      RECT 1011.6000 156.4000 1016.7500 159.4000 ;
      RECT 1003.4500 156.4000 1008.6000 159.4000 ;
      RECT 995.3000 156.4000 1000.4500 159.4000 ;
      RECT 987.1500 156.4000 992.3000 159.4000 ;
      RECT 979.0000 156.4000 984.1500 159.4000 ;
      RECT 970.8500 156.4000 976.0000 159.4000 ;
      RECT 962.7000 156.4000 967.8500 159.4000 ;
      RECT 954.5500 156.4000 959.7000 159.4000 ;
      RECT 946.4000 156.4000 951.5500 159.4000 ;
      RECT 938.2500 156.4000 943.4000 159.4000 ;
      RECT 930.1000 156.4000 935.2500 159.4000 ;
      RECT 921.9500 156.4000 927.1000 159.4000 ;
      RECT 913.8000 156.4000 918.9500 159.4000 ;
      RECT 905.6500 156.4000 910.8000 159.4000 ;
      RECT 897.5000 156.4000 902.6500 159.4000 ;
      RECT 889.3500 156.4000 894.5000 159.4000 ;
      RECT 881.2000 156.4000 886.3500 159.4000 ;
      RECT 873.0500 156.4000 878.2000 159.4000 ;
      RECT 864.9000 156.4000 870.0500 159.4000 ;
      RECT 856.7500 156.4000 861.9000 159.4000 ;
      RECT 848.6000 156.4000 853.7500 159.4000 ;
      RECT 840.4500 156.4000 845.6000 159.4000 ;
      RECT 832.3000 156.4000 837.4500 159.4000 ;
      RECT 824.1500 156.4000 829.3000 159.4000 ;
      RECT 816.0000 156.4000 821.1500 159.4000 ;
      RECT 807.8500 156.4000 813.0000 159.4000 ;
      RECT 799.7000 156.4000 804.8500 159.4000 ;
      RECT 791.5500 156.4000 796.7000 159.4000 ;
      RECT 783.4000 156.4000 788.5500 159.4000 ;
      RECT 775.2500 156.4000 780.4000 159.4000 ;
      RECT 767.1000 156.4000 772.2500 159.4000 ;
      RECT 758.9500 156.4000 764.1000 159.4000 ;
      RECT 750.8000 156.4000 755.9500 159.4000 ;
      RECT 742.6500 156.4000 747.8000 159.4000 ;
      RECT 734.5000 156.4000 739.6500 159.4000 ;
      RECT 726.3500 156.4000 731.5000 159.4000 ;
      RECT 718.2000 156.4000 723.3500 159.4000 ;
      RECT 710.0500 156.4000 715.2000 159.4000 ;
      RECT 701.9000 156.4000 707.0500 159.4000 ;
      RECT 693.7500 156.4000 698.9000 159.4000 ;
      RECT 685.6000 156.4000 690.7500 159.4000 ;
      RECT 677.4500 156.4000 682.6000 159.4000 ;
      RECT 669.3000 156.4000 674.4500 159.4000 ;
      RECT 661.1500 156.4000 666.3000 159.4000 ;
      RECT 653.0000 156.4000 658.1500 159.4000 ;
      RECT 644.8500 156.4000 650.0000 159.4000 ;
      RECT 636.7000 156.4000 641.8500 159.4000 ;
      RECT 628.5500 156.4000 633.7000 159.4000 ;
      RECT 620.4000 156.4000 625.5500 159.4000 ;
      RECT 612.2500 156.4000 617.4000 159.4000 ;
      RECT 604.1000 156.4000 609.2500 159.4000 ;
      RECT 595.9500 156.4000 601.1000 159.4000 ;
      RECT 587.8000 156.4000 592.9500 159.4000 ;
      RECT 579.6500 156.4000 584.8000 159.4000 ;
      RECT 571.5000 156.4000 576.6500 159.4000 ;
      RECT 563.3500 156.4000 568.5000 159.4000 ;
      RECT 555.2000 156.4000 560.3500 159.4000 ;
      RECT 547.0500 156.4000 552.2000 159.4000 ;
      RECT 538.9000 156.4000 544.0500 159.4000 ;
      RECT 530.7500 156.4000 535.9000 159.4000 ;
      RECT 522.6000 156.4000 527.7500 159.4000 ;
      RECT 514.4500 156.4000 519.6000 159.4000 ;
      RECT 506.3000 156.4000 511.4500 159.4000 ;
      RECT 498.1500 156.4000 503.3000 159.4000 ;
      RECT 490.0000 156.4000 495.1500 159.4000 ;
      RECT 481.8500 156.4000 487.0000 159.4000 ;
      RECT 473.7000 156.4000 478.8500 159.4000 ;
      RECT 465.5500 156.4000 470.7000 159.4000 ;
      RECT 457.4000 156.4000 462.5500 159.4000 ;
      RECT 449.2500 156.4000 454.4000 159.4000 ;
      RECT 441.1000 156.4000 446.2500 159.4000 ;
      RECT 432.9500 156.4000 438.1000 159.4000 ;
      RECT 424.8000 156.4000 429.9500 159.4000 ;
      RECT 416.6500 156.4000 421.8000 159.4000 ;
      RECT 396.5000 156.4000 413.6500 159.4000 ;
      RECT 346.5000 156.4000 393.5000 159.4000 ;
      RECT 326.4650 156.4000 343.5000 159.4000 ;
      RECT 317.9500 156.4000 323.4650 159.4000 ;
      RECT 309.4350 156.4000 314.9500 159.4000 ;
      RECT 300.9200 156.4000 306.4350 159.4000 ;
      RECT 292.4050 156.4000 297.9200 159.4000 ;
      RECT 283.8900 156.4000 289.4050 159.4000 ;
      RECT 275.3750 156.4000 280.8900 159.4000 ;
      RECT 266.8600 156.4000 272.3750 159.4000 ;
      RECT 258.3450 156.4000 263.8600 159.4000 ;
      RECT 249.8300 156.4000 255.3450 159.4000 ;
      RECT 241.3150 156.4000 246.8300 159.4000 ;
      RECT 232.8000 156.4000 238.3150 159.4000 ;
      RECT 224.2850 156.4000 229.8000 159.4000 ;
      RECT 215.7700 156.4000 221.2850 159.4000 ;
      RECT 207.2550 156.4000 212.7700 159.4000 ;
      RECT 198.7400 156.4000 204.2550 159.4000 ;
      RECT 190.2250 156.4000 195.7400 159.4000 ;
      RECT 181.7100 156.4000 187.2250 159.4000 ;
      RECT 173.1950 156.4000 178.7100 159.4000 ;
      RECT 164.6800 156.4000 170.1950 159.4000 ;
      RECT 156.1650 156.4000 161.6800 159.4000 ;
      RECT 147.6500 156.4000 153.1650 159.4000 ;
      RECT 139.1350 156.4000 144.6500 159.4000 ;
      RECT 130.6200 156.4000 136.1350 159.4000 ;
      RECT 122.1050 156.4000 127.6200 159.4000 ;
      RECT 113.5900 156.4000 119.1050 159.4000 ;
      RECT 105.0750 156.4000 110.5900 159.4000 ;
      RECT 96.5600 156.4000 102.0750 159.4000 ;
      RECT 88.0450 156.4000 93.5600 159.4000 ;
      RECT 79.5300 156.4000 85.0450 159.4000 ;
      RECT 71.0150 156.4000 76.5300 159.4000 ;
      RECT 62.5000 156.4000 68.0150 159.4000 ;
      RECT 46.5000 156.4000 59.5000 159.4000 ;
      RECT 8.5000 156.4000 43.5000 159.4000 ;
      RECT 0.0000 156.4000 5.5000 159.4000 ;
      RECT 0.0000 154.9000 1120.0000 156.4000 ;
      RECT 1116.6000 154.4000 1120.0000 154.9000 ;
      RECT 0.0000 152.3050 1113.6000 154.9000 ;
      RECT 1118.5000 151.4000 1120.0000 154.4000 ;
      RECT 1114.5000 149.3050 1120.0000 151.4000 ;
      RECT 1076.5000 149.3050 1111.5000 152.3050 ;
      RECT 1060.5000 149.3050 1073.5000 152.3050 ;
      RECT 1052.3500 149.3050 1057.5000 152.3050 ;
      RECT 1044.2000 149.3050 1049.3500 152.3050 ;
      RECT 1036.0500 149.3050 1041.2000 152.3050 ;
      RECT 1027.9000 149.3050 1033.0500 152.3050 ;
      RECT 1019.7500 149.3050 1024.9000 152.3050 ;
      RECT 1011.6000 149.3050 1016.7500 152.3050 ;
      RECT 1003.4500 149.3050 1008.6000 152.3050 ;
      RECT 995.3000 149.3050 1000.4500 152.3050 ;
      RECT 987.1500 149.3050 992.3000 152.3050 ;
      RECT 979.0000 149.3050 984.1500 152.3050 ;
      RECT 970.8500 149.3050 976.0000 152.3050 ;
      RECT 962.7000 149.3050 967.8500 152.3050 ;
      RECT 954.5500 149.3050 959.7000 152.3050 ;
      RECT 946.4000 149.3050 951.5500 152.3050 ;
      RECT 938.2500 149.3050 943.4000 152.3050 ;
      RECT 930.1000 149.3050 935.2500 152.3050 ;
      RECT 921.9500 149.3050 927.1000 152.3050 ;
      RECT 913.8000 149.3050 918.9500 152.3050 ;
      RECT 905.6500 149.3050 910.8000 152.3050 ;
      RECT 897.5000 149.3050 902.6500 152.3050 ;
      RECT 889.3500 149.3050 894.5000 152.3050 ;
      RECT 881.2000 149.3050 886.3500 152.3050 ;
      RECT 873.0500 149.3050 878.2000 152.3050 ;
      RECT 864.9000 149.3050 870.0500 152.3050 ;
      RECT 856.7500 149.3050 861.9000 152.3050 ;
      RECT 848.6000 149.3050 853.7500 152.3050 ;
      RECT 840.4500 149.3050 845.6000 152.3050 ;
      RECT 832.3000 149.3050 837.4500 152.3050 ;
      RECT 824.1500 149.3050 829.3000 152.3050 ;
      RECT 816.0000 149.3050 821.1500 152.3050 ;
      RECT 807.8500 149.3050 813.0000 152.3050 ;
      RECT 799.7000 149.3050 804.8500 152.3050 ;
      RECT 791.5500 149.3050 796.7000 152.3050 ;
      RECT 783.4000 149.3050 788.5500 152.3050 ;
      RECT 775.2500 149.3050 780.4000 152.3050 ;
      RECT 767.1000 149.3050 772.2500 152.3050 ;
      RECT 758.9500 149.3050 764.1000 152.3050 ;
      RECT 750.8000 149.3050 755.9500 152.3050 ;
      RECT 742.6500 149.3050 747.8000 152.3050 ;
      RECT 734.5000 149.3050 739.6500 152.3050 ;
      RECT 726.3500 149.3050 731.5000 152.3050 ;
      RECT 718.2000 149.3050 723.3500 152.3050 ;
      RECT 710.0500 149.3050 715.2000 152.3050 ;
      RECT 701.9000 149.3050 707.0500 152.3050 ;
      RECT 693.7500 149.3050 698.9000 152.3050 ;
      RECT 685.6000 149.3050 690.7500 152.3050 ;
      RECT 677.4500 149.3050 682.6000 152.3050 ;
      RECT 669.3000 149.3050 674.4500 152.3050 ;
      RECT 661.1500 149.3050 666.3000 152.3050 ;
      RECT 653.0000 149.3050 658.1500 152.3050 ;
      RECT 644.8500 149.3050 650.0000 152.3050 ;
      RECT 636.7000 149.3050 641.8500 152.3050 ;
      RECT 628.5500 149.3050 633.7000 152.3050 ;
      RECT 620.4000 149.3050 625.5500 152.3050 ;
      RECT 612.2500 149.3050 617.4000 152.3050 ;
      RECT 604.1000 149.3050 609.2500 152.3050 ;
      RECT 595.9500 149.3050 601.1000 152.3050 ;
      RECT 587.8000 149.3050 592.9500 152.3050 ;
      RECT 579.6500 149.3050 584.8000 152.3050 ;
      RECT 571.5000 149.3050 576.6500 152.3050 ;
      RECT 563.3500 149.3050 568.5000 152.3050 ;
      RECT 555.2000 149.3050 560.3500 152.3050 ;
      RECT 547.0500 149.3050 552.2000 152.3050 ;
      RECT 538.9000 149.3050 544.0500 152.3050 ;
      RECT 530.7500 149.3050 535.9000 152.3050 ;
      RECT 522.6000 149.3050 527.7500 152.3050 ;
      RECT 514.4500 149.3050 519.6000 152.3050 ;
      RECT 506.3000 149.3050 511.4500 152.3050 ;
      RECT 498.1500 149.3050 503.3000 152.3050 ;
      RECT 490.0000 149.3050 495.1500 152.3050 ;
      RECT 481.8500 149.3050 487.0000 152.3050 ;
      RECT 473.7000 149.3050 478.8500 152.3050 ;
      RECT 465.5500 149.3050 470.7000 152.3050 ;
      RECT 457.4000 149.3050 462.5500 152.3050 ;
      RECT 449.2500 149.3050 454.4000 152.3050 ;
      RECT 441.1000 149.3050 446.2500 152.3050 ;
      RECT 432.9500 149.3050 438.1000 152.3050 ;
      RECT 424.8000 149.3050 429.9500 152.3050 ;
      RECT 416.6500 149.3050 421.8000 152.3050 ;
      RECT 396.5000 149.3050 413.6500 152.3050 ;
      RECT 346.5000 149.3050 393.5000 152.3050 ;
      RECT 326.4650 149.3050 343.5000 152.3050 ;
      RECT 317.9500 149.3050 323.4650 152.3050 ;
      RECT 309.4350 149.3050 314.9500 152.3050 ;
      RECT 300.9200 149.3050 306.4350 152.3050 ;
      RECT 292.4050 149.3050 297.9200 152.3050 ;
      RECT 283.8900 149.3050 289.4050 152.3050 ;
      RECT 275.3750 149.3050 280.8900 152.3050 ;
      RECT 266.8600 149.3050 272.3750 152.3050 ;
      RECT 258.3450 149.3050 263.8600 152.3050 ;
      RECT 249.8300 149.3050 255.3450 152.3050 ;
      RECT 241.3150 149.3050 246.8300 152.3050 ;
      RECT 232.8000 149.3050 238.3150 152.3050 ;
      RECT 224.2850 149.3050 229.8000 152.3050 ;
      RECT 215.7700 149.3050 221.2850 152.3050 ;
      RECT 207.2550 149.3050 212.7700 152.3050 ;
      RECT 198.7400 149.3050 204.2550 152.3050 ;
      RECT 190.2250 149.3050 195.7400 152.3050 ;
      RECT 181.7100 149.3050 187.2250 152.3050 ;
      RECT 173.1950 149.3050 178.7100 152.3050 ;
      RECT 164.6800 149.3050 170.1950 152.3050 ;
      RECT 156.1650 149.3050 161.6800 152.3050 ;
      RECT 147.6500 149.3050 153.1650 152.3050 ;
      RECT 139.1350 149.3050 144.6500 152.3050 ;
      RECT 130.6200 149.3050 136.1350 152.3050 ;
      RECT 122.1050 149.3050 127.6200 152.3050 ;
      RECT 113.5900 149.3050 119.1050 152.3050 ;
      RECT 105.0750 149.3050 110.5900 152.3050 ;
      RECT 96.5600 149.3050 102.0750 152.3050 ;
      RECT 88.0450 149.3050 93.5600 152.3050 ;
      RECT 79.5300 149.3050 85.0450 152.3050 ;
      RECT 71.0150 149.3050 76.5300 152.3050 ;
      RECT 62.5000 149.3050 68.0150 152.3050 ;
      RECT 46.5000 149.3050 59.5000 152.3050 ;
      RECT 8.5000 149.3050 43.5000 152.3050 ;
      RECT 0.0000 149.3050 5.5000 152.3050 ;
      RECT 0.0000 147.9000 1120.0000 149.3050 ;
      RECT 1116.6000 147.3050 1120.0000 147.9000 ;
      RECT 0.0000 145.2100 1113.6000 147.9000 ;
      RECT 1118.5000 144.3050 1120.0000 147.3050 ;
      RECT 1114.5000 142.2100 1120.0000 144.3050 ;
      RECT 1076.5000 142.2100 1111.5000 145.2100 ;
      RECT 1060.5000 142.2100 1073.5000 145.2100 ;
      RECT 1052.3500 142.2100 1057.5000 145.2100 ;
      RECT 1044.2000 142.2100 1049.3500 145.2100 ;
      RECT 1036.0500 142.2100 1041.2000 145.2100 ;
      RECT 1027.9000 142.2100 1033.0500 145.2100 ;
      RECT 1019.7500 142.2100 1024.9000 145.2100 ;
      RECT 1011.6000 142.2100 1016.7500 145.2100 ;
      RECT 1003.4500 142.2100 1008.6000 145.2100 ;
      RECT 995.3000 142.2100 1000.4500 145.2100 ;
      RECT 987.1500 142.2100 992.3000 145.2100 ;
      RECT 979.0000 142.2100 984.1500 145.2100 ;
      RECT 970.8500 142.2100 976.0000 145.2100 ;
      RECT 962.7000 142.2100 967.8500 145.2100 ;
      RECT 954.5500 142.2100 959.7000 145.2100 ;
      RECT 946.4000 142.2100 951.5500 145.2100 ;
      RECT 938.2500 142.2100 943.4000 145.2100 ;
      RECT 930.1000 142.2100 935.2500 145.2100 ;
      RECT 921.9500 142.2100 927.1000 145.2100 ;
      RECT 913.8000 142.2100 918.9500 145.2100 ;
      RECT 905.6500 142.2100 910.8000 145.2100 ;
      RECT 897.5000 142.2100 902.6500 145.2100 ;
      RECT 889.3500 142.2100 894.5000 145.2100 ;
      RECT 881.2000 142.2100 886.3500 145.2100 ;
      RECT 873.0500 142.2100 878.2000 145.2100 ;
      RECT 864.9000 142.2100 870.0500 145.2100 ;
      RECT 856.7500 142.2100 861.9000 145.2100 ;
      RECT 848.6000 142.2100 853.7500 145.2100 ;
      RECT 840.4500 142.2100 845.6000 145.2100 ;
      RECT 832.3000 142.2100 837.4500 145.2100 ;
      RECT 824.1500 142.2100 829.3000 145.2100 ;
      RECT 816.0000 142.2100 821.1500 145.2100 ;
      RECT 807.8500 142.2100 813.0000 145.2100 ;
      RECT 799.7000 142.2100 804.8500 145.2100 ;
      RECT 791.5500 142.2100 796.7000 145.2100 ;
      RECT 783.4000 142.2100 788.5500 145.2100 ;
      RECT 775.2500 142.2100 780.4000 145.2100 ;
      RECT 767.1000 142.2100 772.2500 145.2100 ;
      RECT 758.9500 142.2100 764.1000 145.2100 ;
      RECT 750.8000 142.2100 755.9500 145.2100 ;
      RECT 742.6500 142.2100 747.8000 145.2100 ;
      RECT 734.5000 142.2100 739.6500 145.2100 ;
      RECT 726.3500 142.2100 731.5000 145.2100 ;
      RECT 718.2000 142.2100 723.3500 145.2100 ;
      RECT 710.0500 142.2100 715.2000 145.2100 ;
      RECT 701.9000 142.2100 707.0500 145.2100 ;
      RECT 693.7500 142.2100 698.9000 145.2100 ;
      RECT 685.6000 142.2100 690.7500 145.2100 ;
      RECT 677.4500 142.2100 682.6000 145.2100 ;
      RECT 669.3000 142.2100 674.4500 145.2100 ;
      RECT 661.1500 142.2100 666.3000 145.2100 ;
      RECT 653.0000 142.2100 658.1500 145.2100 ;
      RECT 644.8500 142.2100 650.0000 145.2100 ;
      RECT 636.7000 142.2100 641.8500 145.2100 ;
      RECT 628.5500 142.2100 633.7000 145.2100 ;
      RECT 620.4000 142.2100 625.5500 145.2100 ;
      RECT 612.2500 142.2100 617.4000 145.2100 ;
      RECT 604.1000 142.2100 609.2500 145.2100 ;
      RECT 595.9500 142.2100 601.1000 145.2100 ;
      RECT 587.8000 142.2100 592.9500 145.2100 ;
      RECT 579.6500 142.2100 584.8000 145.2100 ;
      RECT 571.5000 142.2100 576.6500 145.2100 ;
      RECT 563.3500 142.2100 568.5000 145.2100 ;
      RECT 555.2000 142.2100 560.3500 145.2100 ;
      RECT 547.0500 142.2100 552.2000 145.2100 ;
      RECT 538.9000 142.2100 544.0500 145.2100 ;
      RECT 530.7500 142.2100 535.9000 145.2100 ;
      RECT 522.6000 142.2100 527.7500 145.2100 ;
      RECT 514.4500 142.2100 519.6000 145.2100 ;
      RECT 506.3000 142.2100 511.4500 145.2100 ;
      RECT 498.1500 142.2100 503.3000 145.2100 ;
      RECT 490.0000 142.2100 495.1500 145.2100 ;
      RECT 481.8500 142.2100 487.0000 145.2100 ;
      RECT 473.7000 142.2100 478.8500 145.2100 ;
      RECT 465.5500 142.2100 470.7000 145.2100 ;
      RECT 457.4000 142.2100 462.5500 145.2100 ;
      RECT 449.2500 142.2100 454.4000 145.2100 ;
      RECT 441.1000 142.2100 446.2500 145.2100 ;
      RECT 432.9500 142.2100 438.1000 145.2100 ;
      RECT 424.8000 142.2100 429.9500 145.2100 ;
      RECT 416.6500 142.2100 421.8000 145.2100 ;
      RECT 396.5000 142.2100 413.6500 145.2100 ;
      RECT 346.5000 142.2100 393.5000 145.2100 ;
      RECT 326.4650 142.2100 343.5000 145.2100 ;
      RECT 317.9500 142.2100 323.4650 145.2100 ;
      RECT 309.4350 142.2100 314.9500 145.2100 ;
      RECT 300.9200 142.2100 306.4350 145.2100 ;
      RECT 292.4050 142.2100 297.9200 145.2100 ;
      RECT 283.8900 142.2100 289.4050 145.2100 ;
      RECT 275.3750 142.2100 280.8900 145.2100 ;
      RECT 266.8600 142.2100 272.3750 145.2100 ;
      RECT 258.3450 142.2100 263.8600 145.2100 ;
      RECT 249.8300 142.2100 255.3450 145.2100 ;
      RECT 241.3150 142.2100 246.8300 145.2100 ;
      RECT 232.8000 142.2100 238.3150 145.2100 ;
      RECT 224.2850 142.2100 229.8000 145.2100 ;
      RECT 215.7700 142.2100 221.2850 145.2100 ;
      RECT 207.2550 142.2100 212.7700 145.2100 ;
      RECT 198.7400 142.2100 204.2550 145.2100 ;
      RECT 190.2250 142.2100 195.7400 145.2100 ;
      RECT 181.7100 142.2100 187.2250 145.2100 ;
      RECT 173.1950 142.2100 178.7100 145.2100 ;
      RECT 164.6800 142.2100 170.1950 145.2100 ;
      RECT 156.1650 142.2100 161.6800 145.2100 ;
      RECT 147.6500 142.2100 153.1650 145.2100 ;
      RECT 139.1350 142.2100 144.6500 145.2100 ;
      RECT 130.6200 142.2100 136.1350 145.2100 ;
      RECT 122.1050 142.2100 127.6200 145.2100 ;
      RECT 113.5900 142.2100 119.1050 145.2100 ;
      RECT 105.0750 142.2100 110.5900 145.2100 ;
      RECT 96.5600 142.2100 102.0750 145.2100 ;
      RECT 88.0450 142.2100 93.5600 145.2100 ;
      RECT 79.5300 142.2100 85.0450 145.2100 ;
      RECT 71.0150 142.2100 76.5300 145.2100 ;
      RECT 62.5000 142.2100 68.0150 145.2100 ;
      RECT 46.5000 142.2100 59.5000 145.2100 ;
      RECT 8.5000 142.2100 43.5000 145.2100 ;
      RECT 0.0000 142.2100 5.5000 145.2100 ;
      RECT 0.0000 140.7000 1120.0000 142.2100 ;
      RECT 1116.6000 140.2100 1120.0000 140.7000 ;
      RECT 0.0000 138.1150 1113.6000 140.7000 ;
      RECT 1118.5000 137.2100 1120.0000 140.2100 ;
      RECT 1114.5000 135.1150 1120.0000 137.2100 ;
      RECT 1076.5000 135.1150 1111.5000 138.1150 ;
      RECT 1060.5000 135.1150 1073.5000 138.1150 ;
      RECT 1052.3500 135.1150 1057.5000 138.1150 ;
      RECT 1044.2000 135.1150 1049.3500 138.1150 ;
      RECT 1036.0500 135.1150 1041.2000 138.1150 ;
      RECT 1027.9000 135.1150 1033.0500 138.1150 ;
      RECT 1019.7500 135.1150 1024.9000 138.1150 ;
      RECT 1011.6000 135.1150 1016.7500 138.1150 ;
      RECT 1003.4500 135.1150 1008.6000 138.1150 ;
      RECT 995.3000 135.1150 1000.4500 138.1150 ;
      RECT 987.1500 135.1150 992.3000 138.1150 ;
      RECT 979.0000 135.1150 984.1500 138.1150 ;
      RECT 970.8500 135.1150 976.0000 138.1150 ;
      RECT 962.7000 135.1150 967.8500 138.1150 ;
      RECT 954.5500 135.1150 959.7000 138.1150 ;
      RECT 946.4000 135.1150 951.5500 138.1150 ;
      RECT 938.2500 135.1150 943.4000 138.1150 ;
      RECT 930.1000 135.1150 935.2500 138.1150 ;
      RECT 921.9500 135.1150 927.1000 138.1150 ;
      RECT 913.8000 135.1150 918.9500 138.1150 ;
      RECT 905.6500 135.1150 910.8000 138.1150 ;
      RECT 897.5000 135.1150 902.6500 138.1150 ;
      RECT 889.3500 135.1150 894.5000 138.1150 ;
      RECT 881.2000 135.1150 886.3500 138.1150 ;
      RECT 873.0500 135.1150 878.2000 138.1150 ;
      RECT 864.9000 135.1150 870.0500 138.1150 ;
      RECT 856.7500 135.1150 861.9000 138.1150 ;
      RECT 848.6000 135.1150 853.7500 138.1150 ;
      RECT 840.4500 135.1150 845.6000 138.1150 ;
      RECT 832.3000 135.1150 837.4500 138.1150 ;
      RECT 824.1500 135.1150 829.3000 138.1150 ;
      RECT 816.0000 135.1150 821.1500 138.1150 ;
      RECT 807.8500 135.1150 813.0000 138.1150 ;
      RECT 799.7000 135.1150 804.8500 138.1150 ;
      RECT 791.5500 135.1150 796.7000 138.1150 ;
      RECT 783.4000 135.1150 788.5500 138.1150 ;
      RECT 775.2500 135.1150 780.4000 138.1150 ;
      RECT 767.1000 135.1150 772.2500 138.1150 ;
      RECT 758.9500 135.1150 764.1000 138.1150 ;
      RECT 750.8000 135.1150 755.9500 138.1150 ;
      RECT 742.6500 135.1150 747.8000 138.1150 ;
      RECT 734.5000 135.1150 739.6500 138.1150 ;
      RECT 726.3500 135.1150 731.5000 138.1150 ;
      RECT 718.2000 135.1150 723.3500 138.1150 ;
      RECT 710.0500 135.1150 715.2000 138.1150 ;
      RECT 701.9000 135.1150 707.0500 138.1150 ;
      RECT 693.7500 135.1150 698.9000 138.1150 ;
      RECT 685.6000 135.1150 690.7500 138.1150 ;
      RECT 677.4500 135.1150 682.6000 138.1150 ;
      RECT 669.3000 135.1150 674.4500 138.1150 ;
      RECT 661.1500 135.1150 666.3000 138.1150 ;
      RECT 653.0000 135.1150 658.1500 138.1150 ;
      RECT 644.8500 135.1150 650.0000 138.1150 ;
      RECT 636.7000 135.1150 641.8500 138.1150 ;
      RECT 628.5500 135.1150 633.7000 138.1150 ;
      RECT 620.4000 135.1150 625.5500 138.1150 ;
      RECT 612.2500 135.1150 617.4000 138.1150 ;
      RECT 604.1000 135.1150 609.2500 138.1150 ;
      RECT 595.9500 135.1150 601.1000 138.1150 ;
      RECT 587.8000 135.1150 592.9500 138.1150 ;
      RECT 579.6500 135.1150 584.8000 138.1150 ;
      RECT 571.5000 135.1150 576.6500 138.1150 ;
      RECT 563.3500 135.1150 568.5000 138.1150 ;
      RECT 555.2000 135.1150 560.3500 138.1150 ;
      RECT 547.0500 135.1150 552.2000 138.1150 ;
      RECT 538.9000 135.1150 544.0500 138.1150 ;
      RECT 530.7500 135.1150 535.9000 138.1150 ;
      RECT 522.6000 135.1150 527.7500 138.1150 ;
      RECT 514.4500 135.1150 519.6000 138.1150 ;
      RECT 506.3000 135.1150 511.4500 138.1150 ;
      RECT 498.1500 135.1150 503.3000 138.1150 ;
      RECT 490.0000 135.1150 495.1500 138.1150 ;
      RECT 481.8500 135.1150 487.0000 138.1150 ;
      RECT 473.7000 135.1150 478.8500 138.1150 ;
      RECT 465.5500 135.1150 470.7000 138.1150 ;
      RECT 457.4000 135.1150 462.5500 138.1150 ;
      RECT 449.2500 135.1150 454.4000 138.1150 ;
      RECT 441.1000 135.1150 446.2500 138.1150 ;
      RECT 432.9500 135.1150 438.1000 138.1150 ;
      RECT 424.8000 135.1150 429.9500 138.1150 ;
      RECT 416.6500 135.1150 421.8000 138.1150 ;
      RECT 396.5000 135.1150 413.6500 138.1150 ;
      RECT 346.5000 135.1150 393.5000 138.1150 ;
      RECT 326.4650 135.1150 343.5000 138.1150 ;
      RECT 317.9500 135.1150 323.4650 138.1150 ;
      RECT 309.4350 135.1150 314.9500 138.1150 ;
      RECT 300.9200 135.1150 306.4350 138.1150 ;
      RECT 292.4050 135.1150 297.9200 138.1150 ;
      RECT 283.8900 135.1150 289.4050 138.1150 ;
      RECT 275.3750 135.1150 280.8900 138.1150 ;
      RECT 266.8600 135.1150 272.3750 138.1150 ;
      RECT 258.3450 135.1150 263.8600 138.1150 ;
      RECT 249.8300 135.1150 255.3450 138.1150 ;
      RECT 241.3150 135.1150 246.8300 138.1150 ;
      RECT 232.8000 135.1150 238.3150 138.1150 ;
      RECT 224.2850 135.1150 229.8000 138.1150 ;
      RECT 215.7700 135.1150 221.2850 138.1150 ;
      RECT 207.2550 135.1150 212.7700 138.1150 ;
      RECT 198.7400 135.1150 204.2550 138.1150 ;
      RECT 190.2250 135.1150 195.7400 138.1150 ;
      RECT 181.7100 135.1150 187.2250 138.1150 ;
      RECT 173.1950 135.1150 178.7100 138.1150 ;
      RECT 164.6800 135.1150 170.1950 138.1150 ;
      RECT 156.1650 135.1150 161.6800 138.1150 ;
      RECT 147.6500 135.1150 153.1650 138.1150 ;
      RECT 139.1350 135.1150 144.6500 138.1150 ;
      RECT 130.6200 135.1150 136.1350 138.1150 ;
      RECT 122.1050 135.1150 127.6200 138.1150 ;
      RECT 113.5900 135.1150 119.1050 138.1150 ;
      RECT 105.0750 135.1150 110.5900 138.1150 ;
      RECT 96.5600 135.1150 102.0750 138.1150 ;
      RECT 88.0450 135.1150 93.5600 138.1150 ;
      RECT 79.5300 135.1150 85.0450 138.1150 ;
      RECT 71.0150 135.1150 76.5300 138.1150 ;
      RECT 62.5000 135.1150 68.0150 138.1150 ;
      RECT 46.5000 135.1150 59.5000 138.1150 ;
      RECT 8.5000 135.1150 43.5000 138.1150 ;
      RECT 0.0000 135.1150 5.5000 138.1150 ;
      RECT 0.0000 133.7000 1120.0000 135.1150 ;
      RECT 1116.6000 133.1150 1120.0000 133.7000 ;
      RECT 0.0000 131.0200 1113.6000 133.7000 ;
      RECT 1118.5000 130.1150 1120.0000 133.1150 ;
      RECT 1114.5000 128.0200 1120.0000 130.1150 ;
      RECT 1076.5000 128.0200 1111.5000 131.0200 ;
      RECT 1060.5000 128.0200 1073.5000 131.0200 ;
      RECT 1052.3500 128.0200 1057.5000 131.0200 ;
      RECT 1044.2000 128.0200 1049.3500 131.0200 ;
      RECT 1036.0500 128.0200 1041.2000 131.0200 ;
      RECT 1027.9000 128.0200 1033.0500 131.0200 ;
      RECT 1019.7500 128.0200 1024.9000 131.0200 ;
      RECT 1011.6000 128.0200 1016.7500 131.0200 ;
      RECT 1003.4500 128.0200 1008.6000 131.0200 ;
      RECT 995.3000 128.0200 1000.4500 131.0200 ;
      RECT 987.1500 128.0200 992.3000 131.0200 ;
      RECT 979.0000 128.0200 984.1500 131.0200 ;
      RECT 970.8500 128.0200 976.0000 131.0200 ;
      RECT 962.7000 128.0200 967.8500 131.0200 ;
      RECT 954.5500 128.0200 959.7000 131.0200 ;
      RECT 946.4000 128.0200 951.5500 131.0200 ;
      RECT 938.2500 128.0200 943.4000 131.0200 ;
      RECT 930.1000 128.0200 935.2500 131.0200 ;
      RECT 921.9500 128.0200 927.1000 131.0200 ;
      RECT 913.8000 128.0200 918.9500 131.0200 ;
      RECT 905.6500 128.0200 910.8000 131.0200 ;
      RECT 897.5000 128.0200 902.6500 131.0200 ;
      RECT 889.3500 128.0200 894.5000 131.0200 ;
      RECT 881.2000 128.0200 886.3500 131.0200 ;
      RECT 873.0500 128.0200 878.2000 131.0200 ;
      RECT 864.9000 128.0200 870.0500 131.0200 ;
      RECT 856.7500 128.0200 861.9000 131.0200 ;
      RECT 848.6000 128.0200 853.7500 131.0200 ;
      RECT 840.4500 128.0200 845.6000 131.0200 ;
      RECT 832.3000 128.0200 837.4500 131.0200 ;
      RECT 824.1500 128.0200 829.3000 131.0200 ;
      RECT 816.0000 128.0200 821.1500 131.0200 ;
      RECT 807.8500 128.0200 813.0000 131.0200 ;
      RECT 799.7000 128.0200 804.8500 131.0200 ;
      RECT 791.5500 128.0200 796.7000 131.0200 ;
      RECT 783.4000 128.0200 788.5500 131.0200 ;
      RECT 775.2500 128.0200 780.4000 131.0200 ;
      RECT 767.1000 128.0200 772.2500 131.0200 ;
      RECT 758.9500 128.0200 764.1000 131.0200 ;
      RECT 750.8000 128.0200 755.9500 131.0200 ;
      RECT 742.6500 128.0200 747.8000 131.0200 ;
      RECT 734.5000 128.0200 739.6500 131.0200 ;
      RECT 726.3500 128.0200 731.5000 131.0200 ;
      RECT 718.2000 128.0200 723.3500 131.0200 ;
      RECT 710.0500 128.0200 715.2000 131.0200 ;
      RECT 701.9000 128.0200 707.0500 131.0200 ;
      RECT 693.7500 128.0200 698.9000 131.0200 ;
      RECT 685.6000 128.0200 690.7500 131.0200 ;
      RECT 677.4500 128.0200 682.6000 131.0200 ;
      RECT 669.3000 128.0200 674.4500 131.0200 ;
      RECT 661.1500 128.0200 666.3000 131.0200 ;
      RECT 653.0000 128.0200 658.1500 131.0200 ;
      RECT 644.8500 128.0200 650.0000 131.0200 ;
      RECT 636.7000 128.0200 641.8500 131.0200 ;
      RECT 628.5500 128.0200 633.7000 131.0200 ;
      RECT 620.4000 128.0200 625.5500 131.0200 ;
      RECT 612.2500 128.0200 617.4000 131.0200 ;
      RECT 604.1000 128.0200 609.2500 131.0200 ;
      RECT 595.9500 128.0200 601.1000 131.0200 ;
      RECT 587.8000 128.0200 592.9500 131.0200 ;
      RECT 579.6500 128.0200 584.8000 131.0200 ;
      RECT 571.5000 128.0200 576.6500 131.0200 ;
      RECT 563.3500 128.0200 568.5000 131.0200 ;
      RECT 555.2000 128.0200 560.3500 131.0200 ;
      RECT 547.0500 128.0200 552.2000 131.0200 ;
      RECT 538.9000 128.0200 544.0500 131.0200 ;
      RECT 530.7500 128.0200 535.9000 131.0200 ;
      RECT 522.6000 128.0200 527.7500 131.0200 ;
      RECT 514.4500 128.0200 519.6000 131.0200 ;
      RECT 506.3000 128.0200 511.4500 131.0200 ;
      RECT 498.1500 128.0200 503.3000 131.0200 ;
      RECT 490.0000 128.0200 495.1500 131.0200 ;
      RECT 481.8500 128.0200 487.0000 131.0200 ;
      RECT 473.7000 128.0200 478.8500 131.0200 ;
      RECT 465.5500 128.0200 470.7000 131.0200 ;
      RECT 457.4000 128.0200 462.5500 131.0200 ;
      RECT 449.2500 128.0200 454.4000 131.0200 ;
      RECT 441.1000 128.0200 446.2500 131.0200 ;
      RECT 432.9500 128.0200 438.1000 131.0200 ;
      RECT 424.8000 128.0200 429.9500 131.0200 ;
      RECT 416.6500 128.0200 421.8000 131.0200 ;
      RECT 396.5000 128.0200 413.6500 131.0200 ;
      RECT 346.5000 128.0200 393.5000 131.0200 ;
      RECT 326.4650 128.0200 343.5000 131.0200 ;
      RECT 317.9500 128.0200 323.4650 131.0200 ;
      RECT 309.4350 128.0200 314.9500 131.0200 ;
      RECT 300.9200 128.0200 306.4350 131.0200 ;
      RECT 292.4050 128.0200 297.9200 131.0200 ;
      RECT 283.8900 128.0200 289.4050 131.0200 ;
      RECT 275.3750 128.0200 280.8900 131.0200 ;
      RECT 266.8600 128.0200 272.3750 131.0200 ;
      RECT 258.3450 128.0200 263.8600 131.0200 ;
      RECT 249.8300 128.0200 255.3450 131.0200 ;
      RECT 241.3150 128.0200 246.8300 131.0200 ;
      RECT 232.8000 128.0200 238.3150 131.0200 ;
      RECT 224.2850 128.0200 229.8000 131.0200 ;
      RECT 215.7700 128.0200 221.2850 131.0200 ;
      RECT 207.2550 128.0200 212.7700 131.0200 ;
      RECT 198.7400 128.0200 204.2550 131.0200 ;
      RECT 190.2250 128.0200 195.7400 131.0200 ;
      RECT 181.7100 128.0200 187.2250 131.0200 ;
      RECT 173.1950 128.0200 178.7100 131.0200 ;
      RECT 164.6800 128.0200 170.1950 131.0200 ;
      RECT 156.1650 128.0200 161.6800 131.0200 ;
      RECT 147.6500 128.0200 153.1650 131.0200 ;
      RECT 139.1350 128.0200 144.6500 131.0200 ;
      RECT 130.6200 128.0200 136.1350 131.0200 ;
      RECT 122.1050 128.0200 127.6200 131.0200 ;
      RECT 113.5900 128.0200 119.1050 131.0200 ;
      RECT 105.0750 128.0200 110.5900 131.0200 ;
      RECT 96.5600 128.0200 102.0750 131.0200 ;
      RECT 88.0450 128.0200 93.5600 131.0200 ;
      RECT 79.5300 128.0200 85.0450 131.0200 ;
      RECT 71.0150 128.0200 76.5300 131.0200 ;
      RECT 62.5000 128.0200 68.0150 131.0200 ;
      RECT 46.5000 128.0200 59.5000 131.0200 ;
      RECT 8.5000 128.0200 43.5000 131.0200 ;
      RECT 0.0000 128.0200 5.5000 131.0200 ;
      RECT 0.0000 126.5000 1120.0000 128.0200 ;
      RECT 1116.6000 126.0200 1120.0000 126.5000 ;
      RECT 0.0000 123.9250 1113.6000 126.5000 ;
      RECT 1118.5000 123.0200 1120.0000 126.0200 ;
      RECT 1114.5000 120.9250 1120.0000 123.0200 ;
      RECT 1076.5000 120.9250 1111.5000 123.9250 ;
      RECT 1060.5000 120.9250 1073.5000 123.9250 ;
      RECT 1052.3500 120.9250 1057.5000 123.9250 ;
      RECT 1044.2000 120.9250 1049.3500 123.9250 ;
      RECT 1036.0500 120.9250 1041.2000 123.9250 ;
      RECT 1027.9000 120.9250 1033.0500 123.9250 ;
      RECT 1019.7500 120.9250 1024.9000 123.9250 ;
      RECT 1011.6000 120.9250 1016.7500 123.9250 ;
      RECT 1003.4500 120.9250 1008.6000 123.9250 ;
      RECT 995.3000 120.9250 1000.4500 123.9250 ;
      RECT 987.1500 120.9250 992.3000 123.9250 ;
      RECT 979.0000 120.9250 984.1500 123.9250 ;
      RECT 970.8500 120.9250 976.0000 123.9250 ;
      RECT 962.7000 120.9250 967.8500 123.9250 ;
      RECT 954.5500 120.9250 959.7000 123.9250 ;
      RECT 946.4000 120.9250 951.5500 123.9250 ;
      RECT 938.2500 120.9250 943.4000 123.9250 ;
      RECT 930.1000 120.9250 935.2500 123.9250 ;
      RECT 921.9500 120.9250 927.1000 123.9250 ;
      RECT 913.8000 120.9250 918.9500 123.9250 ;
      RECT 905.6500 120.9250 910.8000 123.9250 ;
      RECT 897.5000 120.9250 902.6500 123.9250 ;
      RECT 889.3500 120.9250 894.5000 123.9250 ;
      RECT 881.2000 120.9250 886.3500 123.9250 ;
      RECT 873.0500 120.9250 878.2000 123.9250 ;
      RECT 864.9000 120.9250 870.0500 123.9250 ;
      RECT 856.7500 120.9250 861.9000 123.9250 ;
      RECT 848.6000 120.9250 853.7500 123.9250 ;
      RECT 840.4500 120.9250 845.6000 123.9250 ;
      RECT 832.3000 120.9250 837.4500 123.9250 ;
      RECT 824.1500 120.9250 829.3000 123.9250 ;
      RECT 816.0000 120.9250 821.1500 123.9250 ;
      RECT 807.8500 120.9250 813.0000 123.9250 ;
      RECT 799.7000 120.9250 804.8500 123.9250 ;
      RECT 791.5500 120.9250 796.7000 123.9250 ;
      RECT 783.4000 120.9250 788.5500 123.9250 ;
      RECT 775.2500 120.9250 780.4000 123.9250 ;
      RECT 767.1000 120.9250 772.2500 123.9250 ;
      RECT 758.9500 120.9250 764.1000 123.9250 ;
      RECT 750.8000 120.9250 755.9500 123.9250 ;
      RECT 742.6500 120.9250 747.8000 123.9250 ;
      RECT 734.5000 120.9250 739.6500 123.9250 ;
      RECT 726.3500 120.9250 731.5000 123.9250 ;
      RECT 718.2000 120.9250 723.3500 123.9250 ;
      RECT 710.0500 120.9250 715.2000 123.9250 ;
      RECT 701.9000 120.9250 707.0500 123.9250 ;
      RECT 693.7500 120.9250 698.9000 123.9250 ;
      RECT 685.6000 120.9250 690.7500 123.9250 ;
      RECT 677.4500 120.9250 682.6000 123.9250 ;
      RECT 669.3000 120.9250 674.4500 123.9250 ;
      RECT 661.1500 120.9250 666.3000 123.9250 ;
      RECT 653.0000 120.9250 658.1500 123.9250 ;
      RECT 644.8500 120.9250 650.0000 123.9250 ;
      RECT 636.7000 120.9250 641.8500 123.9250 ;
      RECT 628.5500 120.9250 633.7000 123.9250 ;
      RECT 620.4000 120.9250 625.5500 123.9250 ;
      RECT 612.2500 120.9250 617.4000 123.9250 ;
      RECT 604.1000 120.9250 609.2500 123.9250 ;
      RECT 595.9500 120.9250 601.1000 123.9250 ;
      RECT 587.8000 120.9250 592.9500 123.9250 ;
      RECT 579.6500 120.9250 584.8000 123.9250 ;
      RECT 571.5000 120.9250 576.6500 123.9250 ;
      RECT 563.3500 120.9250 568.5000 123.9250 ;
      RECT 555.2000 120.9250 560.3500 123.9250 ;
      RECT 547.0500 120.9250 552.2000 123.9250 ;
      RECT 538.9000 120.9250 544.0500 123.9250 ;
      RECT 530.7500 120.9250 535.9000 123.9250 ;
      RECT 522.6000 120.9250 527.7500 123.9250 ;
      RECT 514.4500 120.9250 519.6000 123.9250 ;
      RECT 506.3000 120.9250 511.4500 123.9250 ;
      RECT 498.1500 120.9250 503.3000 123.9250 ;
      RECT 490.0000 120.9250 495.1500 123.9250 ;
      RECT 481.8500 120.9250 487.0000 123.9250 ;
      RECT 473.7000 120.9250 478.8500 123.9250 ;
      RECT 465.5500 120.9250 470.7000 123.9250 ;
      RECT 457.4000 120.9250 462.5500 123.9250 ;
      RECT 449.2500 120.9250 454.4000 123.9250 ;
      RECT 441.1000 120.9250 446.2500 123.9250 ;
      RECT 432.9500 120.9250 438.1000 123.9250 ;
      RECT 424.8000 120.9250 429.9500 123.9250 ;
      RECT 416.6500 120.9250 421.8000 123.9250 ;
      RECT 396.5000 120.9250 413.6500 123.9250 ;
      RECT 346.5000 120.9250 393.5000 123.9250 ;
      RECT 326.4650 120.9250 343.5000 123.9250 ;
      RECT 317.9500 120.9250 323.4650 123.9250 ;
      RECT 309.4350 120.9250 314.9500 123.9250 ;
      RECT 300.9200 120.9250 306.4350 123.9250 ;
      RECT 292.4050 120.9250 297.9200 123.9250 ;
      RECT 283.8900 120.9250 289.4050 123.9250 ;
      RECT 275.3750 120.9250 280.8900 123.9250 ;
      RECT 266.8600 120.9250 272.3750 123.9250 ;
      RECT 258.3450 120.9250 263.8600 123.9250 ;
      RECT 249.8300 120.9250 255.3450 123.9250 ;
      RECT 241.3150 120.9250 246.8300 123.9250 ;
      RECT 232.8000 120.9250 238.3150 123.9250 ;
      RECT 224.2850 120.9250 229.8000 123.9250 ;
      RECT 215.7700 120.9250 221.2850 123.9250 ;
      RECT 207.2550 120.9250 212.7700 123.9250 ;
      RECT 198.7400 120.9250 204.2550 123.9250 ;
      RECT 190.2250 120.9250 195.7400 123.9250 ;
      RECT 181.7100 120.9250 187.2250 123.9250 ;
      RECT 173.1950 120.9250 178.7100 123.9250 ;
      RECT 164.6800 120.9250 170.1950 123.9250 ;
      RECT 156.1650 120.9250 161.6800 123.9250 ;
      RECT 147.6500 120.9250 153.1650 123.9250 ;
      RECT 139.1350 120.9250 144.6500 123.9250 ;
      RECT 130.6200 120.9250 136.1350 123.9250 ;
      RECT 122.1050 120.9250 127.6200 123.9250 ;
      RECT 113.5900 120.9250 119.1050 123.9250 ;
      RECT 105.0750 120.9250 110.5900 123.9250 ;
      RECT 96.5600 120.9250 102.0750 123.9250 ;
      RECT 88.0450 120.9250 93.5600 123.9250 ;
      RECT 79.5300 120.9250 85.0450 123.9250 ;
      RECT 71.0150 120.9250 76.5300 123.9250 ;
      RECT 62.5000 120.9250 68.0150 123.9250 ;
      RECT 46.5000 120.9250 59.5000 123.9250 ;
      RECT 8.5000 120.9250 43.5000 123.9250 ;
      RECT 0.0000 120.9250 5.5000 123.9250 ;
      RECT 0.0000 119.5000 1120.0000 120.9250 ;
      RECT 1116.6000 118.9250 1120.0000 119.5000 ;
      RECT 0.0000 116.8300 1113.6000 119.5000 ;
      RECT 1118.5000 115.9250 1120.0000 118.9250 ;
      RECT 1114.5000 113.8300 1120.0000 115.9250 ;
      RECT 1076.5000 113.8300 1111.5000 116.8300 ;
      RECT 1060.5000 113.8300 1073.5000 116.8300 ;
      RECT 1052.3500 113.8300 1057.5000 116.8300 ;
      RECT 1044.2000 113.8300 1049.3500 116.8300 ;
      RECT 1036.0500 113.8300 1041.2000 116.8300 ;
      RECT 1027.9000 113.8300 1033.0500 116.8300 ;
      RECT 1019.7500 113.8300 1024.9000 116.8300 ;
      RECT 1011.6000 113.8300 1016.7500 116.8300 ;
      RECT 1003.4500 113.8300 1008.6000 116.8300 ;
      RECT 995.3000 113.8300 1000.4500 116.8300 ;
      RECT 987.1500 113.8300 992.3000 116.8300 ;
      RECT 979.0000 113.8300 984.1500 116.8300 ;
      RECT 970.8500 113.8300 976.0000 116.8300 ;
      RECT 962.7000 113.8300 967.8500 116.8300 ;
      RECT 954.5500 113.8300 959.7000 116.8300 ;
      RECT 946.4000 113.8300 951.5500 116.8300 ;
      RECT 938.2500 113.8300 943.4000 116.8300 ;
      RECT 930.1000 113.8300 935.2500 116.8300 ;
      RECT 921.9500 113.8300 927.1000 116.8300 ;
      RECT 913.8000 113.8300 918.9500 116.8300 ;
      RECT 905.6500 113.8300 910.8000 116.8300 ;
      RECT 897.5000 113.8300 902.6500 116.8300 ;
      RECT 889.3500 113.8300 894.5000 116.8300 ;
      RECT 881.2000 113.8300 886.3500 116.8300 ;
      RECT 873.0500 113.8300 878.2000 116.8300 ;
      RECT 864.9000 113.8300 870.0500 116.8300 ;
      RECT 856.7500 113.8300 861.9000 116.8300 ;
      RECT 848.6000 113.8300 853.7500 116.8300 ;
      RECT 840.4500 113.8300 845.6000 116.8300 ;
      RECT 832.3000 113.8300 837.4500 116.8300 ;
      RECT 824.1500 113.8300 829.3000 116.8300 ;
      RECT 816.0000 113.8300 821.1500 116.8300 ;
      RECT 807.8500 113.8300 813.0000 116.8300 ;
      RECT 799.7000 113.8300 804.8500 116.8300 ;
      RECT 791.5500 113.8300 796.7000 116.8300 ;
      RECT 783.4000 113.8300 788.5500 116.8300 ;
      RECT 775.2500 113.8300 780.4000 116.8300 ;
      RECT 767.1000 113.8300 772.2500 116.8300 ;
      RECT 758.9500 113.8300 764.1000 116.8300 ;
      RECT 750.8000 113.8300 755.9500 116.8300 ;
      RECT 742.6500 113.8300 747.8000 116.8300 ;
      RECT 734.5000 113.8300 739.6500 116.8300 ;
      RECT 726.3500 113.8300 731.5000 116.8300 ;
      RECT 718.2000 113.8300 723.3500 116.8300 ;
      RECT 710.0500 113.8300 715.2000 116.8300 ;
      RECT 701.9000 113.8300 707.0500 116.8300 ;
      RECT 693.7500 113.8300 698.9000 116.8300 ;
      RECT 685.6000 113.8300 690.7500 116.8300 ;
      RECT 677.4500 113.8300 682.6000 116.8300 ;
      RECT 669.3000 113.8300 674.4500 116.8300 ;
      RECT 661.1500 113.8300 666.3000 116.8300 ;
      RECT 653.0000 113.8300 658.1500 116.8300 ;
      RECT 644.8500 113.8300 650.0000 116.8300 ;
      RECT 636.7000 113.8300 641.8500 116.8300 ;
      RECT 628.5500 113.8300 633.7000 116.8300 ;
      RECT 620.4000 113.8300 625.5500 116.8300 ;
      RECT 612.2500 113.8300 617.4000 116.8300 ;
      RECT 604.1000 113.8300 609.2500 116.8300 ;
      RECT 595.9500 113.8300 601.1000 116.8300 ;
      RECT 587.8000 113.8300 592.9500 116.8300 ;
      RECT 579.6500 113.8300 584.8000 116.8300 ;
      RECT 571.5000 113.8300 576.6500 116.8300 ;
      RECT 563.3500 113.8300 568.5000 116.8300 ;
      RECT 555.2000 113.8300 560.3500 116.8300 ;
      RECT 547.0500 113.8300 552.2000 116.8300 ;
      RECT 538.9000 113.8300 544.0500 116.8300 ;
      RECT 530.7500 113.8300 535.9000 116.8300 ;
      RECT 522.6000 113.8300 527.7500 116.8300 ;
      RECT 514.4500 113.8300 519.6000 116.8300 ;
      RECT 506.3000 113.8300 511.4500 116.8300 ;
      RECT 498.1500 113.8300 503.3000 116.8300 ;
      RECT 490.0000 113.8300 495.1500 116.8300 ;
      RECT 481.8500 113.8300 487.0000 116.8300 ;
      RECT 473.7000 113.8300 478.8500 116.8300 ;
      RECT 465.5500 113.8300 470.7000 116.8300 ;
      RECT 457.4000 113.8300 462.5500 116.8300 ;
      RECT 449.2500 113.8300 454.4000 116.8300 ;
      RECT 441.1000 113.8300 446.2500 116.8300 ;
      RECT 432.9500 113.8300 438.1000 116.8300 ;
      RECT 424.8000 113.8300 429.9500 116.8300 ;
      RECT 416.6500 113.8300 421.8000 116.8300 ;
      RECT 396.5000 113.8300 413.6500 116.8300 ;
      RECT 346.5000 113.8300 393.5000 116.8300 ;
      RECT 326.4650 113.8300 343.5000 116.8300 ;
      RECT 317.9500 113.8300 323.4650 116.8300 ;
      RECT 309.4350 113.8300 314.9500 116.8300 ;
      RECT 300.9200 113.8300 306.4350 116.8300 ;
      RECT 292.4050 113.8300 297.9200 116.8300 ;
      RECT 283.8900 113.8300 289.4050 116.8300 ;
      RECT 275.3750 113.8300 280.8900 116.8300 ;
      RECT 266.8600 113.8300 272.3750 116.8300 ;
      RECT 258.3450 113.8300 263.8600 116.8300 ;
      RECT 249.8300 113.8300 255.3450 116.8300 ;
      RECT 241.3150 113.8300 246.8300 116.8300 ;
      RECT 232.8000 113.8300 238.3150 116.8300 ;
      RECT 224.2850 113.8300 229.8000 116.8300 ;
      RECT 215.7700 113.8300 221.2850 116.8300 ;
      RECT 207.2550 113.8300 212.7700 116.8300 ;
      RECT 198.7400 113.8300 204.2550 116.8300 ;
      RECT 190.2250 113.8300 195.7400 116.8300 ;
      RECT 181.7100 113.8300 187.2250 116.8300 ;
      RECT 173.1950 113.8300 178.7100 116.8300 ;
      RECT 164.6800 113.8300 170.1950 116.8300 ;
      RECT 156.1650 113.8300 161.6800 116.8300 ;
      RECT 147.6500 113.8300 153.1650 116.8300 ;
      RECT 139.1350 113.8300 144.6500 116.8300 ;
      RECT 130.6200 113.8300 136.1350 116.8300 ;
      RECT 122.1050 113.8300 127.6200 116.8300 ;
      RECT 113.5900 113.8300 119.1050 116.8300 ;
      RECT 105.0750 113.8300 110.5900 116.8300 ;
      RECT 96.5600 113.8300 102.0750 116.8300 ;
      RECT 88.0450 113.8300 93.5600 116.8300 ;
      RECT 79.5300 113.8300 85.0450 116.8300 ;
      RECT 71.0150 113.8300 76.5300 116.8300 ;
      RECT 62.5000 113.8300 68.0150 116.8300 ;
      RECT 46.5000 113.8300 59.5000 116.8300 ;
      RECT 8.5000 113.8300 43.5000 116.8300 ;
      RECT 0.0000 113.8300 5.5000 116.8300 ;
      RECT 0.0000 112.3000 1120.0000 113.8300 ;
      RECT 1116.6000 111.8300 1120.0000 112.3000 ;
      RECT 0.0000 109.7350 1113.6000 112.3000 ;
      RECT 1118.5000 108.8300 1120.0000 111.8300 ;
      RECT 1114.5000 106.7350 1120.0000 108.8300 ;
      RECT 1076.5000 106.7350 1111.5000 109.7350 ;
      RECT 1060.5000 106.7350 1073.5000 109.7350 ;
      RECT 1052.3500 106.7350 1057.5000 109.7350 ;
      RECT 1044.2000 106.7350 1049.3500 109.7350 ;
      RECT 1036.0500 106.7350 1041.2000 109.7350 ;
      RECT 1027.9000 106.7350 1033.0500 109.7350 ;
      RECT 1019.7500 106.7350 1024.9000 109.7350 ;
      RECT 1011.6000 106.7350 1016.7500 109.7350 ;
      RECT 1003.4500 106.7350 1008.6000 109.7350 ;
      RECT 995.3000 106.7350 1000.4500 109.7350 ;
      RECT 987.1500 106.7350 992.3000 109.7350 ;
      RECT 979.0000 106.7350 984.1500 109.7350 ;
      RECT 970.8500 106.7350 976.0000 109.7350 ;
      RECT 962.7000 106.7350 967.8500 109.7350 ;
      RECT 954.5500 106.7350 959.7000 109.7350 ;
      RECT 946.4000 106.7350 951.5500 109.7350 ;
      RECT 938.2500 106.7350 943.4000 109.7350 ;
      RECT 930.1000 106.7350 935.2500 109.7350 ;
      RECT 921.9500 106.7350 927.1000 109.7350 ;
      RECT 913.8000 106.7350 918.9500 109.7350 ;
      RECT 905.6500 106.7350 910.8000 109.7350 ;
      RECT 897.5000 106.7350 902.6500 109.7350 ;
      RECT 889.3500 106.7350 894.5000 109.7350 ;
      RECT 881.2000 106.7350 886.3500 109.7350 ;
      RECT 873.0500 106.7350 878.2000 109.7350 ;
      RECT 864.9000 106.7350 870.0500 109.7350 ;
      RECT 856.7500 106.7350 861.9000 109.7350 ;
      RECT 848.6000 106.7350 853.7500 109.7350 ;
      RECT 840.4500 106.7350 845.6000 109.7350 ;
      RECT 832.3000 106.7350 837.4500 109.7350 ;
      RECT 824.1500 106.7350 829.3000 109.7350 ;
      RECT 816.0000 106.7350 821.1500 109.7350 ;
      RECT 807.8500 106.7350 813.0000 109.7350 ;
      RECT 799.7000 106.7350 804.8500 109.7350 ;
      RECT 791.5500 106.7350 796.7000 109.7350 ;
      RECT 783.4000 106.7350 788.5500 109.7350 ;
      RECT 775.2500 106.7350 780.4000 109.7350 ;
      RECT 767.1000 106.7350 772.2500 109.7350 ;
      RECT 758.9500 106.7350 764.1000 109.7350 ;
      RECT 750.8000 106.7350 755.9500 109.7350 ;
      RECT 742.6500 106.7350 747.8000 109.7350 ;
      RECT 734.5000 106.7350 739.6500 109.7350 ;
      RECT 726.3500 106.7350 731.5000 109.7350 ;
      RECT 718.2000 106.7350 723.3500 109.7350 ;
      RECT 710.0500 106.7350 715.2000 109.7350 ;
      RECT 701.9000 106.7350 707.0500 109.7350 ;
      RECT 693.7500 106.7350 698.9000 109.7350 ;
      RECT 685.6000 106.7350 690.7500 109.7350 ;
      RECT 677.4500 106.7350 682.6000 109.7350 ;
      RECT 669.3000 106.7350 674.4500 109.7350 ;
      RECT 661.1500 106.7350 666.3000 109.7350 ;
      RECT 653.0000 106.7350 658.1500 109.7350 ;
      RECT 644.8500 106.7350 650.0000 109.7350 ;
      RECT 636.7000 106.7350 641.8500 109.7350 ;
      RECT 628.5500 106.7350 633.7000 109.7350 ;
      RECT 620.4000 106.7350 625.5500 109.7350 ;
      RECT 612.2500 106.7350 617.4000 109.7350 ;
      RECT 604.1000 106.7350 609.2500 109.7350 ;
      RECT 595.9500 106.7350 601.1000 109.7350 ;
      RECT 587.8000 106.7350 592.9500 109.7350 ;
      RECT 579.6500 106.7350 584.8000 109.7350 ;
      RECT 571.5000 106.7350 576.6500 109.7350 ;
      RECT 563.3500 106.7350 568.5000 109.7350 ;
      RECT 555.2000 106.7350 560.3500 109.7350 ;
      RECT 547.0500 106.7350 552.2000 109.7350 ;
      RECT 538.9000 106.7350 544.0500 109.7350 ;
      RECT 530.7500 106.7350 535.9000 109.7350 ;
      RECT 522.6000 106.7350 527.7500 109.7350 ;
      RECT 514.4500 106.7350 519.6000 109.7350 ;
      RECT 506.3000 106.7350 511.4500 109.7350 ;
      RECT 498.1500 106.7350 503.3000 109.7350 ;
      RECT 490.0000 106.7350 495.1500 109.7350 ;
      RECT 481.8500 106.7350 487.0000 109.7350 ;
      RECT 473.7000 106.7350 478.8500 109.7350 ;
      RECT 465.5500 106.7350 470.7000 109.7350 ;
      RECT 457.4000 106.7350 462.5500 109.7350 ;
      RECT 449.2500 106.7350 454.4000 109.7350 ;
      RECT 441.1000 106.7350 446.2500 109.7350 ;
      RECT 432.9500 106.7350 438.1000 109.7350 ;
      RECT 424.8000 106.7350 429.9500 109.7350 ;
      RECT 416.6500 106.7350 421.8000 109.7350 ;
      RECT 396.5000 106.7350 413.6500 109.7350 ;
      RECT 346.5000 106.7350 393.5000 109.7350 ;
      RECT 326.4650 106.7350 343.5000 109.7350 ;
      RECT 317.9500 106.7350 323.4650 109.7350 ;
      RECT 309.4350 106.7350 314.9500 109.7350 ;
      RECT 300.9200 106.7350 306.4350 109.7350 ;
      RECT 292.4050 106.7350 297.9200 109.7350 ;
      RECT 283.8900 106.7350 289.4050 109.7350 ;
      RECT 275.3750 106.7350 280.8900 109.7350 ;
      RECT 266.8600 106.7350 272.3750 109.7350 ;
      RECT 258.3450 106.7350 263.8600 109.7350 ;
      RECT 249.8300 106.7350 255.3450 109.7350 ;
      RECT 241.3150 106.7350 246.8300 109.7350 ;
      RECT 232.8000 106.7350 238.3150 109.7350 ;
      RECT 224.2850 106.7350 229.8000 109.7350 ;
      RECT 215.7700 106.7350 221.2850 109.7350 ;
      RECT 207.2550 106.7350 212.7700 109.7350 ;
      RECT 198.7400 106.7350 204.2550 109.7350 ;
      RECT 190.2250 106.7350 195.7400 109.7350 ;
      RECT 181.7100 106.7350 187.2250 109.7350 ;
      RECT 173.1950 106.7350 178.7100 109.7350 ;
      RECT 164.6800 106.7350 170.1950 109.7350 ;
      RECT 156.1650 106.7350 161.6800 109.7350 ;
      RECT 147.6500 106.7350 153.1650 109.7350 ;
      RECT 139.1350 106.7350 144.6500 109.7350 ;
      RECT 130.6200 106.7350 136.1350 109.7350 ;
      RECT 122.1050 106.7350 127.6200 109.7350 ;
      RECT 113.5900 106.7350 119.1050 109.7350 ;
      RECT 105.0750 106.7350 110.5900 109.7350 ;
      RECT 96.5600 106.7350 102.0750 109.7350 ;
      RECT 88.0450 106.7350 93.5600 109.7350 ;
      RECT 79.5300 106.7350 85.0450 109.7350 ;
      RECT 71.0150 106.7350 76.5300 109.7350 ;
      RECT 62.5000 106.7350 68.0150 109.7350 ;
      RECT 46.5000 106.7350 59.5000 109.7350 ;
      RECT 8.5000 106.7350 43.5000 109.7350 ;
      RECT 0.0000 106.7350 5.5000 109.7350 ;
      RECT 0.0000 105.3000 1120.0000 106.7350 ;
      RECT 1116.6000 104.7350 1120.0000 105.3000 ;
      RECT 0.0000 102.6400 1113.6000 105.3000 ;
      RECT 1118.5000 101.7350 1120.0000 104.7350 ;
      RECT 1114.5000 99.6400 1120.0000 101.7350 ;
      RECT 1076.5000 99.6400 1111.5000 102.6400 ;
      RECT 1060.5000 99.6400 1073.5000 102.6400 ;
      RECT 1052.3500 99.6400 1057.5000 102.6400 ;
      RECT 1044.2000 99.6400 1049.3500 102.6400 ;
      RECT 1036.0500 99.6400 1041.2000 102.6400 ;
      RECT 1027.9000 99.6400 1033.0500 102.6400 ;
      RECT 1019.7500 99.6400 1024.9000 102.6400 ;
      RECT 1011.6000 99.6400 1016.7500 102.6400 ;
      RECT 1003.4500 99.6400 1008.6000 102.6400 ;
      RECT 995.3000 99.6400 1000.4500 102.6400 ;
      RECT 987.1500 99.6400 992.3000 102.6400 ;
      RECT 979.0000 99.6400 984.1500 102.6400 ;
      RECT 970.8500 99.6400 976.0000 102.6400 ;
      RECT 962.7000 99.6400 967.8500 102.6400 ;
      RECT 954.5500 99.6400 959.7000 102.6400 ;
      RECT 946.4000 99.6400 951.5500 102.6400 ;
      RECT 938.2500 99.6400 943.4000 102.6400 ;
      RECT 930.1000 99.6400 935.2500 102.6400 ;
      RECT 921.9500 99.6400 927.1000 102.6400 ;
      RECT 913.8000 99.6400 918.9500 102.6400 ;
      RECT 905.6500 99.6400 910.8000 102.6400 ;
      RECT 897.5000 99.6400 902.6500 102.6400 ;
      RECT 889.3500 99.6400 894.5000 102.6400 ;
      RECT 881.2000 99.6400 886.3500 102.6400 ;
      RECT 873.0500 99.6400 878.2000 102.6400 ;
      RECT 864.9000 99.6400 870.0500 102.6400 ;
      RECT 856.7500 99.6400 861.9000 102.6400 ;
      RECT 848.6000 99.6400 853.7500 102.6400 ;
      RECT 840.4500 99.6400 845.6000 102.6400 ;
      RECT 832.3000 99.6400 837.4500 102.6400 ;
      RECT 824.1500 99.6400 829.3000 102.6400 ;
      RECT 816.0000 99.6400 821.1500 102.6400 ;
      RECT 807.8500 99.6400 813.0000 102.6400 ;
      RECT 799.7000 99.6400 804.8500 102.6400 ;
      RECT 791.5500 99.6400 796.7000 102.6400 ;
      RECT 783.4000 99.6400 788.5500 102.6400 ;
      RECT 775.2500 99.6400 780.4000 102.6400 ;
      RECT 767.1000 99.6400 772.2500 102.6400 ;
      RECT 758.9500 99.6400 764.1000 102.6400 ;
      RECT 750.8000 99.6400 755.9500 102.6400 ;
      RECT 742.6500 99.6400 747.8000 102.6400 ;
      RECT 734.5000 99.6400 739.6500 102.6400 ;
      RECT 726.3500 99.6400 731.5000 102.6400 ;
      RECT 718.2000 99.6400 723.3500 102.6400 ;
      RECT 710.0500 99.6400 715.2000 102.6400 ;
      RECT 701.9000 99.6400 707.0500 102.6400 ;
      RECT 693.7500 99.6400 698.9000 102.6400 ;
      RECT 685.6000 99.6400 690.7500 102.6400 ;
      RECT 677.4500 99.6400 682.6000 102.6400 ;
      RECT 669.3000 99.6400 674.4500 102.6400 ;
      RECT 661.1500 99.6400 666.3000 102.6400 ;
      RECT 653.0000 99.6400 658.1500 102.6400 ;
      RECT 644.8500 99.6400 650.0000 102.6400 ;
      RECT 636.7000 99.6400 641.8500 102.6400 ;
      RECT 628.5500 99.6400 633.7000 102.6400 ;
      RECT 620.4000 99.6400 625.5500 102.6400 ;
      RECT 612.2500 99.6400 617.4000 102.6400 ;
      RECT 604.1000 99.6400 609.2500 102.6400 ;
      RECT 595.9500 99.6400 601.1000 102.6400 ;
      RECT 587.8000 99.6400 592.9500 102.6400 ;
      RECT 579.6500 99.6400 584.8000 102.6400 ;
      RECT 571.5000 99.6400 576.6500 102.6400 ;
      RECT 563.3500 99.6400 568.5000 102.6400 ;
      RECT 555.2000 99.6400 560.3500 102.6400 ;
      RECT 547.0500 99.6400 552.2000 102.6400 ;
      RECT 538.9000 99.6400 544.0500 102.6400 ;
      RECT 530.7500 99.6400 535.9000 102.6400 ;
      RECT 522.6000 99.6400 527.7500 102.6400 ;
      RECT 514.4500 99.6400 519.6000 102.6400 ;
      RECT 506.3000 99.6400 511.4500 102.6400 ;
      RECT 498.1500 99.6400 503.3000 102.6400 ;
      RECT 490.0000 99.6400 495.1500 102.6400 ;
      RECT 481.8500 99.6400 487.0000 102.6400 ;
      RECT 473.7000 99.6400 478.8500 102.6400 ;
      RECT 465.5500 99.6400 470.7000 102.6400 ;
      RECT 457.4000 99.6400 462.5500 102.6400 ;
      RECT 449.2500 99.6400 454.4000 102.6400 ;
      RECT 441.1000 99.6400 446.2500 102.6400 ;
      RECT 432.9500 99.6400 438.1000 102.6400 ;
      RECT 424.8000 99.6400 429.9500 102.6400 ;
      RECT 416.6500 99.6400 421.8000 102.6400 ;
      RECT 396.5000 99.6400 413.6500 102.6400 ;
      RECT 346.5000 99.6400 393.5000 102.6400 ;
      RECT 326.4650 99.6400 343.5000 102.6400 ;
      RECT 317.9500 99.6400 323.4650 102.6400 ;
      RECT 309.4350 99.6400 314.9500 102.6400 ;
      RECT 300.9200 99.6400 306.4350 102.6400 ;
      RECT 292.4050 99.6400 297.9200 102.6400 ;
      RECT 283.8900 99.6400 289.4050 102.6400 ;
      RECT 275.3750 99.6400 280.8900 102.6400 ;
      RECT 266.8600 99.6400 272.3750 102.6400 ;
      RECT 258.3450 99.6400 263.8600 102.6400 ;
      RECT 249.8300 99.6400 255.3450 102.6400 ;
      RECT 241.3150 99.6400 246.8300 102.6400 ;
      RECT 232.8000 99.6400 238.3150 102.6400 ;
      RECT 224.2850 99.6400 229.8000 102.6400 ;
      RECT 215.7700 99.6400 221.2850 102.6400 ;
      RECT 207.2550 99.6400 212.7700 102.6400 ;
      RECT 198.7400 99.6400 204.2550 102.6400 ;
      RECT 190.2250 99.6400 195.7400 102.6400 ;
      RECT 181.7100 99.6400 187.2250 102.6400 ;
      RECT 173.1950 99.6400 178.7100 102.6400 ;
      RECT 164.6800 99.6400 170.1950 102.6400 ;
      RECT 156.1650 99.6400 161.6800 102.6400 ;
      RECT 147.6500 99.6400 153.1650 102.6400 ;
      RECT 139.1350 99.6400 144.6500 102.6400 ;
      RECT 130.6200 99.6400 136.1350 102.6400 ;
      RECT 122.1050 99.6400 127.6200 102.6400 ;
      RECT 113.5900 99.6400 119.1050 102.6400 ;
      RECT 105.0750 99.6400 110.5900 102.6400 ;
      RECT 96.5600 99.6400 102.0750 102.6400 ;
      RECT 88.0450 99.6400 93.5600 102.6400 ;
      RECT 79.5300 99.6400 85.0450 102.6400 ;
      RECT 71.0150 99.6400 76.5300 102.6400 ;
      RECT 62.5000 99.6400 68.0150 102.6400 ;
      RECT 46.5000 99.6400 59.5000 102.6400 ;
      RECT 8.5000 99.6400 43.5000 102.6400 ;
      RECT 0.0000 99.6400 5.5000 102.6400 ;
      RECT 0.0000 98.1000 1120.0000 99.6400 ;
      RECT 1116.6000 97.6400 1120.0000 98.1000 ;
      RECT 0.0000 95.5450 1113.6000 98.1000 ;
      RECT 1118.5000 94.6400 1120.0000 97.6400 ;
      RECT 1114.5000 92.5450 1120.0000 94.6400 ;
      RECT 1076.5000 92.5450 1111.5000 95.5450 ;
      RECT 1060.5000 92.5450 1073.5000 95.5450 ;
      RECT 1052.3500 92.5450 1057.5000 95.5450 ;
      RECT 1044.2000 92.5450 1049.3500 95.5450 ;
      RECT 1036.0500 92.5450 1041.2000 95.5450 ;
      RECT 1027.9000 92.5450 1033.0500 95.5450 ;
      RECT 1019.7500 92.5450 1024.9000 95.5450 ;
      RECT 1011.6000 92.5450 1016.7500 95.5450 ;
      RECT 1003.4500 92.5450 1008.6000 95.5450 ;
      RECT 995.3000 92.5450 1000.4500 95.5450 ;
      RECT 987.1500 92.5450 992.3000 95.5450 ;
      RECT 979.0000 92.5450 984.1500 95.5450 ;
      RECT 970.8500 92.5450 976.0000 95.5450 ;
      RECT 962.7000 92.5450 967.8500 95.5450 ;
      RECT 954.5500 92.5450 959.7000 95.5450 ;
      RECT 946.4000 92.5450 951.5500 95.5450 ;
      RECT 938.2500 92.5450 943.4000 95.5450 ;
      RECT 930.1000 92.5450 935.2500 95.5450 ;
      RECT 921.9500 92.5450 927.1000 95.5450 ;
      RECT 913.8000 92.5450 918.9500 95.5450 ;
      RECT 905.6500 92.5450 910.8000 95.5450 ;
      RECT 897.5000 92.5450 902.6500 95.5450 ;
      RECT 889.3500 92.5450 894.5000 95.5450 ;
      RECT 881.2000 92.5450 886.3500 95.5450 ;
      RECT 873.0500 92.5450 878.2000 95.5450 ;
      RECT 864.9000 92.5450 870.0500 95.5450 ;
      RECT 856.7500 92.5450 861.9000 95.5450 ;
      RECT 848.6000 92.5450 853.7500 95.5450 ;
      RECT 840.4500 92.5450 845.6000 95.5450 ;
      RECT 832.3000 92.5450 837.4500 95.5450 ;
      RECT 824.1500 92.5450 829.3000 95.5450 ;
      RECT 816.0000 92.5450 821.1500 95.5450 ;
      RECT 807.8500 92.5450 813.0000 95.5450 ;
      RECT 799.7000 92.5450 804.8500 95.5450 ;
      RECT 791.5500 92.5450 796.7000 95.5450 ;
      RECT 783.4000 92.5450 788.5500 95.5450 ;
      RECT 775.2500 92.5450 780.4000 95.5450 ;
      RECT 767.1000 92.5450 772.2500 95.5450 ;
      RECT 758.9500 92.5450 764.1000 95.5450 ;
      RECT 750.8000 92.5450 755.9500 95.5450 ;
      RECT 742.6500 92.5450 747.8000 95.5450 ;
      RECT 734.5000 92.5450 739.6500 95.5450 ;
      RECT 726.3500 92.5450 731.5000 95.5450 ;
      RECT 718.2000 92.5450 723.3500 95.5450 ;
      RECT 710.0500 92.5450 715.2000 95.5450 ;
      RECT 701.9000 92.5450 707.0500 95.5450 ;
      RECT 693.7500 92.5450 698.9000 95.5450 ;
      RECT 685.6000 92.5450 690.7500 95.5450 ;
      RECT 677.4500 92.5450 682.6000 95.5450 ;
      RECT 669.3000 92.5450 674.4500 95.5450 ;
      RECT 661.1500 92.5450 666.3000 95.5450 ;
      RECT 653.0000 92.5450 658.1500 95.5450 ;
      RECT 644.8500 92.5450 650.0000 95.5450 ;
      RECT 636.7000 92.5450 641.8500 95.5450 ;
      RECT 628.5500 92.5450 633.7000 95.5450 ;
      RECT 620.4000 92.5450 625.5500 95.5450 ;
      RECT 612.2500 92.5450 617.4000 95.5450 ;
      RECT 604.1000 92.5450 609.2500 95.5450 ;
      RECT 595.9500 92.5450 601.1000 95.5450 ;
      RECT 587.8000 92.5450 592.9500 95.5450 ;
      RECT 579.6500 92.5450 584.8000 95.5450 ;
      RECT 571.5000 92.5450 576.6500 95.5450 ;
      RECT 563.3500 92.5450 568.5000 95.5450 ;
      RECT 555.2000 92.5450 560.3500 95.5450 ;
      RECT 547.0500 92.5450 552.2000 95.5450 ;
      RECT 538.9000 92.5450 544.0500 95.5450 ;
      RECT 530.7500 92.5450 535.9000 95.5450 ;
      RECT 522.6000 92.5450 527.7500 95.5450 ;
      RECT 514.4500 92.5450 519.6000 95.5450 ;
      RECT 506.3000 92.5450 511.4500 95.5450 ;
      RECT 498.1500 92.5450 503.3000 95.5450 ;
      RECT 490.0000 92.5450 495.1500 95.5450 ;
      RECT 481.8500 92.5450 487.0000 95.5450 ;
      RECT 473.7000 92.5450 478.8500 95.5450 ;
      RECT 465.5500 92.5450 470.7000 95.5450 ;
      RECT 457.4000 92.5450 462.5500 95.5450 ;
      RECT 449.2500 92.5450 454.4000 95.5450 ;
      RECT 441.1000 92.5450 446.2500 95.5450 ;
      RECT 432.9500 92.5450 438.1000 95.5450 ;
      RECT 424.8000 92.5450 429.9500 95.5450 ;
      RECT 416.6500 92.5450 421.8000 95.5450 ;
      RECT 396.5000 92.5450 413.6500 95.5450 ;
      RECT 346.5000 92.5450 393.5000 95.5450 ;
      RECT 326.4650 92.5450 343.5000 95.5450 ;
      RECT 317.9500 92.5450 323.4650 95.5450 ;
      RECT 309.4350 92.5450 314.9500 95.5450 ;
      RECT 300.9200 92.5450 306.4350 95.5450 ;
      RECT 292.4050 92.5450 297.9200 95.5450 ;
      RECT 283.8900 92.5450 289.4050 95.5450 ;
      RECT 275.3750 92.5450 280.8900 95.5450 ;
      RECT 266.8600 92.5450 272.3750 95.5450 ;
      RECT 258.3450 92.5450 263.8600 95.5450 ;
      RECT 249.8300 92.5450 255.3450 95.5450 ;
      RECT 241.3150 92.5450 246.8300 95.5450 ;
      RECT 232.8000 92.5450 238.3150 95.5450 ;
      RECT 224.2850 92.5450 229.8000 95.5450 ;
      RECT 215.7700 92.5450 221.2850 95.5450 ;
      RECT 207.2550 92.5450 212.7700 95.5450 ;
      RECT 198.7400 92.5450 204.2550 95.5450 ;
      RECT 190.2250 92.5450 195.7400 95.5450 ;
      RECT 181.7100 92.5450 187.2250 95.5450 ;
      RECT 173.1950 92.5450 178.7100 95.5450 ;
      RECT 164.6800 92.5450 170.1950 95.5450 ;
      RECT 156.1650 92.5450 161.6800 95.5450 ;
      RECT 147.6500 92.5450 153.1650 95.5450 ;
      RECT 139.1350 92.5450 144.6500 95.5450 ;
      RECT 130.6200 92.5450 136.1350 95.5450 ;
      RECT 122.1050 92.5450 127.6200 95.5450 ;
      RECT 113.5900 92.5450 119.1050 95.5450 ;
      RECT 105.0750 92.5450 110.5900 95.5450 ;
      RECT 96.5600 92.5450 102.0750 95.5450 ;
      RECT 88.0450 92.5450 93.5600 95.5450 ;
      RECT 79.5300 92.5450 85.0450 95.5450 ;
      RECT 71.0150 92.5450 76.5300 95.5450 ;
      RECT 62.5000 92.5450 68.0150 95.5450 ;
      RECT 46.5000 92.5450 59.5000 95.5450 ;
      RECT 8.5000 92.5450 43.5000 95.5450 ;
      RECT 0.0000 92.5450 5.5000 95.5450 ;
      RECT 0.0000 91.1000 1120.0000 92.5450 ;
      RECT 1116.6000 90.5450 1120.0000 91.1000 ;
      RECT 0.0000 88.4500 1113.6000 91.1000 ;
      RECT 1118.5000 87.5450 1120.0000 90.5450 ;
      RECT 1114.5000 85.4500 1120.0000 87.5450 ;
      RECT 1076.5000 85.4500 1111.5000 88.4500 ;
      RECT 1060.5000 85.4500 1073.5000 88.4500 ;
      RECT 1052.3500 85.4500 1057.5000 88.4500 ;
      RECT 1044.2000 85.4500 1049.3500 88.4500 ;
      RECT 1036.0500 85.4500 1041.2000 88.4500 ;
      RECT 1027.9000 85.4500 1033.0500 88.4500 ;
      RECT 1019.7500 85.4500 1024.9000 88.4500 ;
      RECT 1011.6000 85.4500 1016.7500 88.4500 ;
      RECT 1003.4500 85.4500 1008.6000 88.4500 ;
      RECT 995.3000 85.4500 1000.4500 88.4500 ;
      RECT 987.1500 85.4500 992.3000 88.4500 ;
      RECT 979.0000 85.4500 984.1500 88.4500 ;
      RECT 970.8500 85.4500 976.0000 88.4500 ;
      RECT 962.7000 85.4500 967.8500 88.4500 ;
      RECT 954.5500 85.4500 959.7000 88.4500 ;
      RECT 946.4000 85.4500 951.5500 88.4500 ;
      RECT 938.2500 85.4500 943.4000 88.4500 ;
      RECT 930.1000 85.4500 935.2500 88.4500 ;
      RECT 921.9500 85.4500 927.1000 88.4500 ;
      RECT 913.8000 85.4500 918.9500 88.4500 ;
      RECT 905.6500 85.4500 910.8000 88.4500 ;
      RECT 897.5000 85.4500 902.6500 88.4500 ;
      RECT 889.3500 85.4500 894.5000 88.4500 ;
      RECT 881.2000 85.4500 886.3500 88.4500 ;
      RECT 873.0500 85.4500 878.2000 88.4500 ;
      RECT 864.9000 85.4500 870.0500 88.4500 ;
      RECT 856.7500 85.4500 861.9000 88.4500 ;
      RECT 848.6000 85.4500 853.7500 88.4500 ;
      RECT 840.4500 85.4500 845.6000 88.4500 ;
      RECT 832.3000 85.4500 837.4500 88.4500 ;
      RECT 824.1500 85.4500 829.3000 88.4500 ;
      RECT 816.0000 85.4500 821.1500 88.4500 ;
      RECT 807.8500 85.4500 813.0000 88.4500 ;
      RECT 799.7000 85.4500 804.8500 88.4500 ;
      RECT 791.5500 85.4500 796.7000 88.4500 ;
      RECT 783.4000 85.4500 788.5500 88.4500 ;
      RECT 775.2500 85.4500 780.4000 88.4500 ;
      RECT 767.1000 85.4500 772.2500 88.4500 ;
      RECT 758.9500 85.4500 764.1000 88.4500 ;
      RECT 750.8000 85.4500 755.9500 88.4500 ;
      RECT 742.6500 85.4500 747.8000 88.4500 ;
      RECT 734.5000 85.4500 739.6500 88.4500 ;
      RECT 726.3500 85.4500 731.5000 88.4500 ;
      RECT 718.2000 85.4500 723.3500 88.4500 ;
      RECT 710.0500 85.4500 715.2000 88.4500 ;
      RECT 701.9000 85.4500 707.0500 88.4500 ;
      RECT 693.7500 85.4500 698.9000 88.4500 ;
      RECT 685.6000 85.4500 690.7500 88.4500 ;
      RECT 677.4500 85.4500 682.6000 88.4500 ;
      RECT 669.3000 85.4500 674.4500 88.4500 ;
      RECT 661.1500 85.4500 666.3000 88.4500 ;
      RECT 653.0000 85.4500 658.1500 88.4500 ;
      RECT 644.8500 85.4500 650.0000 88.4500 ;
      RECT 636.7000 85.4500 641.8500 88.4500 ;
      RECT 628.5500 85.4500 633.7000 88.4500 ;
      RECT 620.4000 85.4500 625.5500 88.4500 ;
      RECT 612.2500 85.4500 617.4000 88.4500 ;
      RECT 604.1000 85.4500 609.2500 88.4500 ;
      RECT 595.9500 85.4500 601.1000 88.4500 ;
      RECT 587.8000 85.4500 592.9500 88.4500 ;
      RECT 579.6500 85.4500 584.8000 88.4500 ;
      RECT 571.5000 85.4500 576.6500 88.4500 ;
      RECT 563.3500 85.4500 568.5000 88.4500 ;
      RECT 555.2000 85.4500 560.3500 88.4500 ;
      RECT 547.0500 85.4500 552.2000 88.4500 ;
      RECT 538.9000 85.4500 544.0500 88.4500 ;
      RECT 530.7500 85.4500 535.9000 88.4500 ;
      RECT 522.6000 85.4500 527.7500 88.4500 ;
      RECT 514.4500 85.4500 519.6000 88.4500 ;
      RECT 506.3000 85.4500 511.4500 88.4500 ;
      RECT 498.1500 85.4500 503.3000 88.4500 ;
      RECT 490.0000 85.4500 495.1500 88.4500 ;
      RECT 481.8500 85.4500 487.0000 88.4500 ;
      RECT 473.7000 85.4500 478.8500 88.4500 ;
      RECT 465.5500 85.4500 470.7000 88.4500 ;
      RECT 457.4000 85.4500 462.5500 88.4500 ;
      RECT 449.2500 85.4500 454.4000 88.4500 ;
      RECT 441.1000 85.4500 446.2500 88.4500 ;
      RECT 432.9500 85.4500 438.1000 88.4500 ;
      RECT 424.8000 85.4500 429.9500 88.4500 ;
      RECT 416.6500 85.4500 421.8000 88.4500 ;
      RECT 396.5000 85.4500 413.6500 88.4500 ;
      RECT 346.5000 85.4500 393.5000 88.4500 ;
      RECT 326.4650 85.4500 343.5000 88.4500 ;
      RECT 317.9500 85.4500 323.4650 88.4500 ;
      RECT 309.4350 85.4500 314.9500 88.4500 ;
      RECT 300.9200 85.4500 306.4350 88.4500 ;
      RECT 292.4050 85.4500 297.9200 88.4500 ;
      RECT 283.8900 85.4500 289.4050 88.4500 ;
      RECT 275.3750 85.4500 280.8900 88.4500 ;
      RECT 266.8600 85.4500 272.3750 88.4500 ;
      RECT 258.3450 85.4500 263.8600 88.4500 ;
      RECT 249.8300 85.4500 255.3450 88.4500 ;
      RECT 241.3150 85.4500 246.8300 88.4500 ;
      RECT 232.8000 85.4500 238.3150 88.4500 ;
      RECT 224.2850 85.4500 229.8000 88.4500 ;
      RECT 215.7700 85.4500 221.2850 88.4500 ;
      RECT 207.2550 85.4500 212.7700 88.4500 ;
      RECT 198.7400 85.4500 204.2550 88.4500 ;
      RECT 190.2250 85.4500 195.7400 88.4500 ;
      RECT 181.7100 85.4500 187.2250 88.4500 ;
      RECT 173.1950 85.4500 178.7100 88.4500 ;
      RECT 164.6800 85.4500 170.1950 88.4500 ;
      RECT 156.1650 85.4500 161.6800 88.4500 ;
      RECT 147.6500 85.4500 153.1650 88.4500 ;
      RECT 139.1350 85.4500 144.6500 88.4500 ;
      RECT 130.6200 85.4500 136.1350 88.4500 ;
      RECT 122.1050 85.4500 127.6200 88.4500 ;
      RECT 113.5900 85.4500 119.1050 88.4500 ;
      RECT 105.0750 85.4500 110.5900 88.4500 ;
      RECT 96.5600 85.4500 102.0750 88.4500 ;
      RECT 88.0450 85.4500 93.5600 88.4500 ;
      RECT 79.5300 85.4500 85.0450 88.4500 ;
      RECT 71.0150 85.4500 76.5300 88.4500 ;
      RECT 62.5000 85.4500 68.0150 88.4500 ;
      RECT 46.5000 85.4500 59.5000 88.4500 ;
      RECT 8.5000 85.4500 43.5000 88.4500 ;
      RECT 0.0000 85.4500 5.5000 88.4500 ;
      RECT 0.0000 83.9000 1120.0000 85.4500 ;
      RECT 1116.6000 83.4500 1120.0000 83.9000 ;
      RECT 0.0000 81.3550 1113.6000 83.9000 ;
      RECT 1118.5000 80.4500 1120.0000 83.4500 ;
      RECT 1114.5000 78.3550 1120.0000 80.4500 ;
      RECT 1076.5000 78.3550 1111.5000 81.3550 ;
      RECT 1060.5000 78.3550 1073.5000 81.3550 ;
      RECT 1052.3500 78.3550 1057.5000 81.3550 ;
      RECT 1044.2000 78.3550 1049.3500 81.3550 ;
      RECT 1036.0500 78.3550 1041.2000 81.3550 ;
      RECT 1027.9000 78.3550 1033.0500 81.3550 ;
      RECT 1019.7500 78.3550 1024.9000 81.3550 ;
      RECT 1011.6000 78.3550 1016.7500 81.3550 ;
      RECT 1003.4500 78.3550 1008.6000 81.3550 ;
      RECT 995.3000 78.3550 1000.4500 81.3550 ;
      RECT 987.1500 78.3550 992.3000 81.3550 ;
      RECT 979.0000 78.3550 984.1500 81.3550 ;
      RECT 970.8500 78.3550 976.0000 81.3550 ;
      RECT 962.7000 78.3550 967.8500 81.3550 ;
      RECT 954.5500 78.3550 959.7000 81.3550 ;
      RECT 946.4000 78.3550 951.5500 81.3550 ;
      RECT 938.2500 78.3550 943.4000 81.3550 ;
      RECT 930.1000 78.3550 935.2500 81.3550 ;
      RECT 921.9500 78.3550 927.1000 81.3550 ;
      RECT 913.8000 78.3550 918.9500 81.3550 ;
      RECT 905.6500 78.3550 910.8000 81.3550 ;
      RECT 897.5000 78.3550 902.6500 81.3550 ;
      RECT 889.3500 78.3550 894.5000 81.3550 ;
      RECT 881.2000 78.3550 886.3500 81.3550 ;
      RECT 873.0500 78.3550 878.2000 81.3550 ;
      RECT 864.9000 78.3550 870.0500 81.3550 ;
      RECT 856.7500 78.3550 861.9000 81.3550 ;
      RECT 848.6000 78.3550 853.7500 81.3550 ;
      RECT 840.4500 78.3550 845.6000 81.3550 ;
      RECT 832.3000 78.3550 837.4500 81.3550 ;
      RECT 824.1500 78.3550 829.3000 81.3550 ;
      RECT 816.0000 78.3550 821.1500 81.3550 ;
      RECT 807.8500 78.3550 813.0000 81.3550 ;
      RECT 799.7000 78.3550 804.8500 81.3550 ;
      RECT 791.5500 78.3550 796.7000 81.3550 ;
      RECT 783.4000 78.3550 788.5500 81.3550 ;
      RECT 775.2500 78.3550 780.4000 81.3550 ;
      RECT 767.1000 78.3550 772.2500 81.3550 ;
      RECT 758.9500 78.3550 764.1000 81.3550 ;
      RECT 750.8000 78.3550 755.9500 81.3550 ;
      RECT 742.6500 78.3550 747.8000 81.3550 ;
      RECT 734.5000 78.3550 739.6500 81.3550 ;
      RECT 726.3500 78.3550 731.5000 81.3550 ;
      RECT 718.2000 78.3550 723.3500 81.3550 ;
      RECT 710.0500 78.3550 715.2000 81.3550 ;
      RECT 701.9000 78.3550 707.0500 81.3550 ;
      RECT 693.7500 78.3550 698.9000 81.3550 ;
      RECT 685.6000 78.3550 690.7500 81.3550 ;
      RECT 677.4500 78.3550 682.6000 81.3550 ;
      RECT 669.3000 78.3550 674.4500 81.3550 ;
      RECT 661.1500 78.3550 666.3000 81.3550 ;
      RECT 653.0000 78.3550 658.1500 81.3550 ;
      RECT 644.8500 78.3550 650.0000 81.3550 ;
      RECT 636.7000 78.3550 641.8500 81.3550 ;
      RECT 628.5500 78.3550 633.7000 81.3550 ;
      RECT 620.4000 78.3550 625.5500 81.3550 ;
      RECT 612.2500 78.3550 617.4000 81.3550 ;
      RECT 604.1000 78.3550 609.2500 81.3550 ;
      RECT 595.9500 78.3550 601.1000 81.3550 ;
      RECT 587.8000 78.3550 592.9500 81.3550 ;
      RECT 579.6500 78.3550 584.8000 81.3550 ;
      RECT 571.5000 78.3550 576.6500 81.3550 ;
      RECT 563.3500 78.3550 568.5000 81.3550 ;
      RECT 555.2000 78.3550 560.3500 81.3550 ;
      RECT 547.0500 78.3550 552.2000 81.3550 ;
      RECT 538.9000 78.3550 544.0500 81.3550 ;
      RECT 530.7500 78.3550 535.9000 81.3550 ;
      RECT 522.6000 78.3550 527.7500 81.3550 ;
      RECT 514.4500 78.3550 519.6000 81.3550 ;
      RECT 506.3000 78.3550 511.4500 81.3550 ;
      RECT 498.1500 78.3550 503.3000 81.3550 ;
      RECT 490.0000 78.3550 495.1500 81.3550 ;
      RECT 481.8500 78.3550 487.0000 81.3550 ;
      RECT 473.7000 78.3550 478.8500 81.3550 ;
      RECT 465.5500 78.3550 470.7000 81.3550 ;
      RECT 457.4000 78.3550 462.5500 81.3550 ;
      RECT 449.2500 78.3550 454.4000 81.3550 ;
      RECT 441.1000 78.3550 446.2500 81.3550 ;
      RECT 432.9500 78.3550 438.1000 81.3550 ;
      RECT 424.8000 78.3550 429.9500 81.3550 ;
      RECT 416.6500 78.3550 421.8000 81.3550 ;
      RECT 396.5000 78.3550 413.6500 81.3550 ;
      RECT 346.5000 78.3550 393.5000 81.3550 ;
      RECT 326.4650 78.3550 343.5000 81.3550 ;
      RECT 317.9500 78.3550 323.4650 81.3550 ;
      RECT 309.4350 78.3550 314.9500 81.3550 ;
      RECT 300.9200 78.3550 306.4350 81.3550 ;
      RECT 292.4050 78.3550 297.9200 81.3550 ;
      RECT 283.8900 78.3550 289.4050 81.3550 ;
      RECT 275.3750 78.3550 280.8900 81.3550 ;
      RECT 266.8600 78.3550 272.3750 81.3550 ;
      RECT 258.3450 78.3550 263.8600 81.3550 ;
      RECT 249.8300 78.3550 255.3450 81.3550 ;
      RECT 241.3150 78.3550 246.8300 81.3550 ;
      RECT 232.8000 78.3550 238.3150 81.3550 ;
      RECT 224.2850 78.3550 229.8000 81.3550 ;
      RECT 215.7700 78.3550 221.2850 81.3550 ;
      RECT 207.2550 78.3550 212.7700 81.3550 ;
      RECT 198.7400 78.3550 204.2550 81.3550 ;
      RECT 190.2250 78.3550 195.7400 81.3550 ;
      RECT 181.7100 78.3550 187.2250 81.3550 ;
      RECT 173.1950 78.3550 178.7100 81.3550 ;
      RECT 164.6800 78.3550 170.1950 81.3550 ;
      RECT 156.1650 78.3550 161.6800 81.3550 ;
      RECT 147.6500 78.3550 153.1650 81.3550 ;
      RECT 139.1350 78.3550 144.6500 81.3550 ;
      RECT 130.6200 78.3550 136.1350 81.3550 ;
      RECT 122.1050 78.3550 127.6200 81.3550 ;
      RECT 113.5900 78.3550 119.1050 81.3550 ;
      RECT 105.0750 78.3550 110.5900 81.3550 ;
      RECT 96.5600 78.3550 102.0750 81.3550 ;
      RECT 88.0450 78.3550 93.5600 81.3550 ;
      RECT 79.5300 78.3550 85.0450 81.3550 ;
      RECT 71.0150 78.3550 76.5300 81.3550 ;
      RECT 62.5000 78.3550 68.0150 81.3550 ;
      RECT 46.5000 78.3550 59.5000 81.3550 ;
      RECT 8.5000 78.3550 43.5000 81.3550 ;
      RECT 0.0000 78.3550 5.5000 81.3550 ;
      RECT 0.0000 76.9000 1120.0000 78.3550 ;
      RECT 1116.6000 76.3550 1120.0000 76.9000 ;
      RECT 0.0000 74.2600 1113.6000 76.9000 ;
      RECT 1118.5000 73.3550 1120.0000 76.3550 ;
      RECT 1114.5000 71.2600 1120.0000 73.3550 ;
      RECT 1076.5000 71.2600 1111.5000 74.2600 ;
      RECT 1060.5000 71.2600 1073.5000 74.2600 ;
      RECT 1052.3500 71.2600 1057.5000 74.2600 ;
      RECT 1044.2000 71.2600 1049.3500 74.2600 ;
      RECT 1036.0500 71.2600 1041.2000 74.2600 ;
      RECT 1027.9000 71.2600 1033.0500 74.2600 ;
      RECT 1019.7500 71.2600 1024.9000 74.2600 ;
      RECT 1011.6000 71.2600 1016.7500 74.2600 ;
      RECT 1003.4500 71.2600 1008.6000 74.2600 ;
      RECT 995.3000 71.2600 1000.4500 74.2600 ;
      RECT 987.1500 71.2600 992.3000 74.2600 ;
      RECT 979.0000 71.2600 984.1500 74.2600 ;
      RECT 970.8500 71.2600 976.0000 74.2600 ;
      RECT 962.7000 71.2600 967.8500 74.2600 ;
      RECT 954.5500 71.2600 959.7000 74.2600 ;
      RECT 946.4000 71.2600 951.5500 74.2600 ;
      RECT 938.2500 71.2600 943.4000 74.2600 ;
      RECT 930.1000 71.2600 935.2500 74.2600 ;
      RECT 921.9500 71.2600 927.1000 74.2600 ;
      RECT 913.8000 71.2600 918.9500 74.2600 ;
      RECT 905.6500 71.2600 910.8000 74.2600 ;
      RECT 897.5000 71.2600 902.6500 74.2600 ;
      RECT 889.3500 71.2600 894.5000 74.2600 ;
      RECT 881.2000 71.2600 886.3500 74.2600 ;
      RECT 873.0500 71.2600 878.2000 74.2600 ;
      RECT 864.9000 71.2600 870.0500 74.2600 ;
      RECT 856.7500 71.2600 861.9000 74.2600 ;
      RECT 848.6000 71.2600 853.7500 74.2600 ;
      RECT 840.4500 71.2600 845.6000 74.2600 ;
      RECT 832.3000 71.2600 837.4500 74.2600 ;
      RECT 824.1500 71.2600 829.3000 74.2600 ;
      RECT 816.0000 71.2600 821.1500 74.2600 ;
      RECT 807.8500 71.2600 813.0000 74.2600 ;
      RECT 799.7000 71.2600 804.8500 74.2600 ;
      RECT 791.5500 71.2600 796.7000 74.2600 ;
      RECT 783.4000 71.2600 788.5500 74.2600 ;
      RECT 775.2500 71.2600 780.4000 74.2600 ;
      RECT 767.1000 71.2600 772.2500 74.2600 ;
      RECT 758.9500 71.2600 764.1000 74.2600 ;
      RECT 750.8000 71.2600 755.9500 74.2600 ;
      RECT 742.6500 71.2600 747.8000 74.2600 ;
      RECT 734.5000 71.2600 739.6500 74.2600 ;
      RECT 726.3500 71.2600 731.5000 74.2600 ;
      RECT 718.2000 71.2600 723.3500 74.2600 ;
      RECT 710.0500 71.2600 715.2000 74.2600 ;
      RECT 701.9000 71.2600 707.0500 74.2600 ;
      RECT 693.7500 71.2600 698.9000 74.2600 ;
      RECT 685.6000 71.2600 690.7500 74.2600 ;
      RECT 677.4500 71.2600 682.6000 74.2600 ;
      RECT 669.3000 71.2600 674.4500 74.2600 ;
      RECT 661.1500 71.2600 666.3000 74.2600 ;
      RECT 653.0000 71.2600 658.1500 74.2600 ;
      RECT 644.8500 71.2600 650.0000 74.2600 ;
      RECT 636.7000 71.2600 641.8500 74.2600 ;
      RECT 628.5500 71.2600 633.7000 74.2600 ;
      RECT 620.4000 71.2600 625.5500 74.2600 ;
      RECT 612.2500 71.2600 617.4000 74.2600 ;
      RECT 604.1000 71.2600 609.2500 74.2600 ;
      RECT 595.9500 71.2600 601.1000 74.2600 ;
      RECT 587.8000 71.2600 592.9500 74.2600 ;
      RECT 579.6500 71.2600 584.8000 74.2600 ;
      RECT 571.5000 71.2600 576.6500 74.2600 ;
      RECT 563.3500 71.2600 568.5000 74.2600 ;
      RECT 555.2000 71.2600 560.3500 74.2600 ;
      RECT 547.0500 71.2600 552.2000 74.2600 ;
      RECT 538.9000 71.2600 544.0500 74.2600 ;
      RECT 530.7500 71.2600 535.9000 74.2600 ;
      RECT 522.6000 71.2600 527.7500 74.2600 ;
      RECT 514.4500 71.2600 519.6000 74.2600 ;
      RECT 506.3000 71.2600 511.4500 74.2600 ;
      RECT 498.1500 71.2600 503.3000 74.2600 ;
      RECT 490.0000 71.2600 495.1500 74.2600 ;
      RECT 481.8500 71.2600 487.0000 74.2600 ;
      RECT 473.7000 71.2600 478.8500 74.2600 ;
      RECT 465.5500 71.2600 470.7000 74.2600 ;
      RECT 457.4000 71.2600 462.5500 74.2600 ;
      RECT 449.2500 71.2600 454.4000 74.2600 ;
      RECT 441.1000 71.2600 446.2500 74.2600 ;
      RECT 432.9500 71.2600 438.1000 74.2600 ;
      RECT 424.8000 71.2600 429.9500 74.2600 ;
      RECT 416.6500 71.2600 421.8000 74.2600 ;
      RECT 396.5000 71.2600 413.6500 74.2600 ;
      RECT 346.5000 71.2600 393.5000 74.2600 ;
      RECT 326.4650 71.2600 343.5000 74.2600 ;
      RECT 317.9500 71.2600 323.4650 74.2600 ;
      RECT 309.4350 71.2600 314.9500 74.2600 ;
      RECT 300.9200 71.2600 306.4350 74.2600 ;
      RECT 292.4050 71.2600 297.9200 74.2600 ;
      RECT 283.8900 71.2600 289.4050 74.2600 ;
      RECT 275.3750 71.2600 280.8900 74.2600 ;
      RECT 266.8600 71.2600 272.3750 74.2600 ;
      RECT 258.3450 71.2600 263.8600 74.2600 ;
      RECT 249.8300 71.2600 255.3450 74.2600 ;
      RECT 241.3150 71.2600 246.8300 74.2600 ;
      RECT 232.8000 71.2600 238.3150 74.2600 ;
      RECT 224.2850 71.2600 229.8000 74.2600 ;
      RECT 215.7700 71.2600 221.2850 74.2600 ;
      RECT 207.2550 71.2600 212.7700 74.2600 ;
      RECT 198.7400 71.2600 204.2550 74.2600 ;
      RECT 190.2250 71.2600 195.7400 74.2600 ;
      RECT 181.7100 71.2600 187.2250 74.2600 ;
      RECT 173.1950 71.2600 178.7100 74.2600 ;
      RECT 164.6800 71.2600 170.1950 74.2600 ;
      RECT 156.1650 71.2600 161.6800 74.2600 ;
      RECT 147.6500 71.2600 153.1650 74.2600 ;
      RECT 139.1350 71.2600 144.6500 74.2600 ;
      RECT 130.6200 71.2600 136.1350 74.2600 ;
      RECT 122.1050 71.2600 127.6200 74.2600 ;
      RECT 113.5900 71.2600 119.1050 74.2600 ;
      RECT 105.0750 71.2600 110.5900 74.2600 ;
      RECT 96.5600 71.2600 102.0750 74.2600 ;
      RECT 88.0450 71.2600 93.5600 74.2600 ;
      RECT 79.5300 71.2600 85.0450 74.2600 ;
      RECT 71.0150 71.2600 76.5300 74.2600 ;
      RECT 62.5000 71.2600 68.0150 74.2600 ;
      RECT 46.5000 71.2600 59.5000 74.2600 ;
      RECT 8.5000 71.2600 43.5000 74.2600 ;
      RECT 0.0000 71.2600 5.5000 74.2600 ;
      RECT 0.0000 69.7000 1120.0000 71.2600 ;
      RECT 1116.6000 69.2600 1120.0000 69.7000 ;
      RECT 0.0000 67.1650 1113.6000 69.7000 ;
      RECT 1118.5000 66.2600 1120.0000 69.2600 ;
      RECT 1114.5000 64.1650 1120.0000 66.2600 ;
      RECT 1076.5000 64.1650 1111.5000 67.1650 ;
      RECT 1060.5000 64.1650 1073.5000 67.1650 ;
      RECT 1052.3500 64.1650 1057.5000 67.1650 ;
      RECT 1044.2000 64.1650 1049.3500 67.1650 ;
      RECT 1036.0500 64.1650 1041.2000 67.1650 ;
      RECT 1027.9000 64.1650 1033.0500 67.1650 ;
      RECT 1019.7500 64.1650 1024.9000 67.1650 ;
      RECT 1011.6000 64.1650 1016.7500 67.1650 ;
      RECT 1003.4500 64.1650 1008.6000 67.1650 ;
      RECT 995.3000 64.1650 1000.4500 67.1650 ;
      RECT 987.1500 64.1650 992.3000 67.1650 ;
      RECT 979.0000 64.1650 984.1500 67.1650 ;
      RECT 970.8500 64.1650 976.0000 67.1650 ;
      RECT 962.7000 64.1650 967.8500 67.1650 ;
      RECT 954.5500 64.1650 959.7000 67.1650 ;
      RECT 946.4000 64.1650 951.5500 67.1650 ;
      RECT 938.2500 64.1650 943.4000 67.1650 ;
      RECT 930.1000 64.1650 935.2500 67.1650 ;
      RECT 921.9500 64.1650 927.1000 67.1650 ;
      RECT 913.8000 64.1650 918.9500 67.1650 ;
      RECT 905.6500 64.1650 910.8000 67.1650 ;
      RECT 897.5000 64.1650 902.6500 67.1650 ;
      RECT 889.3500 64.1650 894.5000 67.1650 ;
      RECT 881.2000 64.1650 886.3500 67.1650 ;
      RECT 873.0500 64.1650 878.2000 67.1650 ;
      RECT 864.9000 64.1650 870.0500 67.1650 ;
      RECT 856.7500 64.1650 861.9000 67.1650 ;
      RECT 848.6000 64.1650 853.7500 67.1650 ;
      RECT 840.4500 64.1650 845.6000 67.1650 ;
      RECT 832.3000 64.1650 837.4500 67.1650 ;
      RECT 824.1500 64.1650 829.3000 67.1650 ;
      RECT 816.0000 64.1650 821.1500 67.1650 ;
      RECT 807.8500 64.1650 813.0000 67.1650 ;
      RECT 799.7000 64.1650 804.8500 67.1650 ;
      RECT 791.5500 64.1650 796.7000 67.1650 ;
      RECT 783.4000 64.1650 788.5500 67.1650 ;
      RECT 775.2500 64.1650 780.4000 67.1650 ;
      RECT 767.1000 64.1650 772.2500 67.1650 ;
      RECT 758.9500 64.1650 764.1000 67.1650 ;
      RECT 750.8000 64.1650 755.9500 67.1650 ;
      RECT 742.6500 64.1650 747.8000 67.1650 ;
      RECT 734.5000 64.1650 739.6500 67.1650 ;
      RECT 726.3500 64.1650 731.5000 67.1650 ;
      RECT 718.2000 64.1650 723.3500 67.1650 ;
      RECT 710.0500 64.1650 715.2000 67.1650 ;
      RECT 701.9000 64.1650 707.0500 67.1650 ;
      RECT 693.7500 64.1650 698.9000 67.1650 ;
      RECT 685.6000 64.1650 690.7500 67.1650 ;
      RECT 677.4500 64.1650 682.6000 67.1650 ;
      RECT 669.3000 64.1650 674.4500 67.1650 ;
      RECT 661.1500 64.1650 666.3000 67.1650 ;
      RECT 653.0000 64.1650 658.1500 67.1650 ;
      RECT 644.8500 64.1650 650.0000 67.1650 ;
      RECT 636.7000 64.1650 641.8500 67.1650 ;
      RECT 628.5500 64.1650 633.7000 67.1650 ;
      RECT 620.4000 64.1650 625.5500 67.1650 ;
      RECT 612.2500 64.1650 617.4000 67.1650 ;
      RECT 604.1000 64.1650 609.2500 67.1650 ;
      RECT 595.9500 64.1650 601.1000 67.1650 ;
      RECT 587.8000 64.1650 592.9500 67.1650 ;
      RECT 579.6500 64.1650 584.8000 67.1650 ;
      RECT 571.5000 64.1650 576.6500 67.1650 ;
      RECT 563.3500 64.1650 568.5000 67.1650 ;
      RECT 555.2000 64.1650 560.3500 67.1650 ;
      RECT 547.0500 64.1650 552.2000 67.1650 ;
      RECT 538.9000 64.1650 544.0500 67.1650 ;
      RECT 530.7500 64.1650 535.9000 67.1650 ;
      RECT 522.6000 64.1650 527.7500 67.1650 ;
      RECT 514.4500 64.1650 519.6000 67.1650 ;
      RECT 506.3000 64.1650 511.4500 67.1650 ;
      RECT 498.1500 64.1650 503.3000 67.1650 ;
      RECT 490.0000 64.1650 495.1500 67.1650 ;
      RECT 481.8500 64.1650 487.0000 67.1650 ;
      RECT 473.7000 64.1650 478.8500 67.1650 ;
      RECT 465.5500 64.1650 470.7000 67.1650 ;
      RECT 457.4000 64.1650 462.5500 67.1650 ;
      RECT 449.2500 64.1650 454.4000 67.1650 ;
      RECT 441.1000 64.1650 446.2500 67.1650 ;
      RECT 432.9500 64.1650 438.1000 67.1650 ;
      RECT 424.8000 64.1650 429.9500 67.1650 ;
      RECT 416.6500 64.1650 421.8000 67.1650 ;
      RECT 396.5000 64.1650 413.6500 67.1650 ;
      RECT 346.5000 64.1650 393.5000 67.1650 ;
      RECT 326.4650 64.1650 343.5000 67.1650 ;
      RECT 317.9500 64.1650 323.4650 67.1650 ;
      RECT 309.4350 64.1650 314.9500 67.1650 ;
      RECT 300.9200 64.1650 306.4350 67.1650 ;
      RECT 292.4050 64.1650 297.9200 67.1650 ;
      RECT 283.8900 64.1650 289.4050 67.1650 ;
      RECT 275.3750 64.1650 280.8900 67.1650 ;
      RECT 266.8600 64.1650 272.3750 67.1650 ;
      RECT 258.3450 64.1650 263.8600 67.1650 ;
      RECT 249.8300 64.1650 255.3450 67.1650 ;
      RECT 241.3150 64.1650 246.8300 67.1650 ;
      RECT 232.8000 64.1650 238.3150 67.1650 ;
      RECT 224.2850 64.1650 229.8000 67.1650 ;
      RECT 215.7700 64.1650 221.2850 67.1650 ;
      RECT 207.2550 64.1650 212.7700 67.1650 ;
      RECT 198.7400 64.1650 204.2550 67.1650 ;
      RECT 190.2250 64.1650 195.7400 67.1650 ;
      RECT 181.7100 64.1650 187.2250 67.1650 ;
      RECT 173.1950 64.1650 178.7100 67.1650 ;
      RECT 164.6800 64.1650 170.1950 67.1650 ;
      RECT 156.1650 64.1650 161.6800 67.1650 ;
      RECT 147.6500 64.1650 153.1650 67.1650 ;
      RECT 139.1350 64.1650 144.6500 67.1650 ;
      RECT 130.6200 64.1650 136.1350 67.1650 ;
      RECT 122.1050 64.1650 127.6200 67.1650 ;
      RECT 113.5900 64.1650 119.1050 67.1650 ;
      RECT 105.0750 64.1650 110.5900 67.1650 ;
      RECT 96.5600 64.1650 102.0750 67.1650 ;
      RECT 88.0450 64.1650 93.5600 67.1650 ;
      RECT 79.5300 64.1650 85.0450 67.1650 ;
      RECT 71.0150 64.1650 76.5300 67.1650 ;
      RECT 62.5000 64.1650 68.0150 67.1650 ;
      RECT 46.5000 64.1650 59.5000 67.1650 ;
      RECT 8.5000 64.1650 43.5000 67.1650 ;
      RECT 0.0000 64.1650 5.5000 67.1650 ;
      RECT 0.0000 62.7000 1120.0000 64.1650 ;
      RECT 0.0000 62.5000 1113.6000 62.7000 ;
      RECT 62.5000 62.3350 1113.6000 62.5000 ;
      RECT 1116.6000 62.1650 1120.0000 62.7000 ;
      RECT 109.0750 60.0700 1113.6000 62.3350 ;
      RECT 0.0000 60.0700 59.5000 62.5000 ;
      RECT 109.0750 59.5700 343.5000 60.0700 ;
      RECT 62.5000 59.5700 106.0750 62.3350 ;
      RECT 62.5000 59.5000 343.5000 59.5700 ;
      RECT 46.5000 59.5000 59.5000 60.0700 ;
      RECT 1118.5000 59.1650 1120.0000 62.1650 ;
      RECT 1114.5000 57.0700 1120.0000 59.1650 ;
      RECT 1076.5000 57.0700 1111.5000 60.0700 ;
      RECT 396.5000 57.0700 1073.5000 60.0700 ;
      RECT 346.5000 57.0700 393.5000 60.0700 ;
      RECT 46.5000 57.0700 343.5000 59.5000 ;
      RECT 8.5000 57.0700 43.5000 60.0700 ;
      RECT 0.0000 57.0700 5.5000 60.0700 ;
      RECT 0.0000 55.5000 1120.0000 57.0700 ;
      RECT 1116.6000 55.0700 1120.0000 55.5000 ;
      RECT 0.0000 52.9750 1113.6000 55.5000 ;
      RECT 1118.5000 52.0700 1120.0000 55.0700 ;
      RECT 1114.5000 49.9750 1120.0000 52.0700 ;
      RECT 1076.5000 49.9750 1111.5000 52.9750 ;
      RECT 396.5000 49.9750 1073.5000 52.9750 ;
      RECT 346.5000 49.9750 393.5000 52.9750 ;
      RECT 46.5000 49.9750 343.5000 52.9750 ;
      RECT 8.5000 49.9750 43.5000 52.9750 ;
      RECT 0.0000 49.9750 5.5000 52.9750 ;
      RECT 0.0000 49.5000 1120.0000 49.9750 ;
      RECT 1116.6000 47.9750 1120.0000 49.5000 ;
      RECT 109.0750 46.5000 1113.6000 49.5000 ;
      RECT 0.0000 46.5000 106.0750 49.5000 ;
      RECT 0.0000 45.8800 1113.6000 46.5000 ;
      RECT 1118.5000 44.9750 1120.0000 47.9750 ;
      RECT 1076.5000 43.5000 1111.5000 45.8800 ;
      RECT 396.5000 43.5000 1073.5000 45.8800 ;
      RECT 346.5000 43.5000 393.5000 45.8800 ;
      RECT 46.5000 43.5000 343.5000 45.8800 ;
      RECT 8.5000 43.5000 43.5000 45.8800 ;
      RECT 1114.5000 42.8800 1120.0000 44.9750 ;
      RECT 8.5000 42.8800 1111.5000 43.5000 ;
      RECT 0.0000 42.8800 5.5000 45.8800 ;
      RECT 0.0000 40.8800 1120.0000 42.8800 ;
      RECT 0.0000 38.7850 1114.0000 40.8800 ;
      RECT 1118.5000 37.8800 1120.0000 40.8800 ;
      RECT 8.5000 35.7850 1111.5000 38.7850 ;
      RECT 0.0000 35.7850 5.5000 38.7850 ;
      RECT 1117.0000 33.7850 1120.0000 37.8800 ;
      RECT 0.0000 31.6900 1114.0000 35.7850 ;
      RECT 1118.5000 30.7850 1120.0000 33.7850 ;
      RECT 8.5000 28.6900 1111.5000 31.6900 ;
      RECT 0.0000 28.6900 5.5000 31.6900 ;
      RECT 1117.0000 26.6900 1120.0000 30.7850 ;
      RECT 0.0000 24.5950 1114.0000 28.6900 ;
      RECT 1118.5000 23.6900 1120.0000 26.6900 ;
      RECT 8.5000 21.5950 1111.5000 24.5950 ;
      RECT 0.0000 21.5950 5.5000 24.5950 ;
      RECT 1117.0000 19.5950 1120.0000 23.6900 ;
      RECT 0.0000 17.5000 1114.0000 21.5950 ;
      RECT 1118.5000 16.5950 1120.0000 19.5950 ;
      RECT 8.5000 14.5000 1111.5000 17.5000 ;
      RECT 0.0000 14.5000 5.5000 17.5000 ;
      RECT 1117.0000 12.5000 1120.0000 16.5950 ;
      RECT 0.0000 12.5000 1114.0000 14.5000 ;
      RECT 1118.5000 9.5000 1120.0000 12.5000 ;
      RECT 4.5000 9.5000 1114.0000 12.5000 ;
      RECT 0.0000 9.5000 1.5000 12.5000 ;
      RECT 1117.0000 1.5000 1120.0000 9.5000 ;
      RECT 0.0000 1.5000 1114.0000 9.5000 ;
      RECT 0.0000 0.0000 1120.0000 1.5000 ;
  END
END core

END LIBRARY
