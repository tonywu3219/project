##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 20:48:30 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 1420.0000 BY 2820.0000 ;
  FOREIGN fullchip 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1369.7500 0.5200 1369.8500 ;
    END
  END clk
  PIN mem_in_core0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1407.7500 0.5200 1407.8500 ;
    END
  END mem_in_core0[63]
  PIN mem_in_core0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1403.7500 0.5200 1403.8500 ;
    END
  END mem_in_core0[62]
  PIN mem_in_core0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1399.7500 0.5200 1399.8500 ;
    END
  END mem_in_core0[61]
  PIN mem_in_core0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1395.7500 0.5200 1395.8500 ;
    END
  END mem_in_core0[60]
  PIN mem_in_core0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1391.7500 0.5200 1391.8500 ;
    END
  END mem_in_core0[59]
  PIN mem_in_core0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1387.7500 0.5200 1387.8500 ;
    END
  END mem_in_core0[58]
  PIN mem_in_core0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1383.7500 0.5200 1383.8500 ;
    END
  END mem_in_core0[57]
  PIN mem_in_core0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1379.7500 0.5200 1379.8500 ;
    END
  END mem_in_core0[56]
  PIN mem_in_core0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1375.7500 0.5200 1375.8500 ;
    END
  END mem_in_core0[55]
  PIN mem_in_core0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1371.7500 0.5200 1371.8500 ;
    END
  END mem_in_core0[54]
  PIN mem_in_core0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1367.7500 0.5200 1367.8500 ;
    END
  END mem_in_core0[53]
  PIN mem_in_core0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1363.7500 0.5200 1363.8500 ;
    END
  END mem_in_core0[52]
  PIN mem_in_core0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1359.7500 0.5200 1359.8500 ;
    END
  END mem_in_core0[51]
  PIN mem_in_core0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1355.7500 0.5200 1355.8500 ;
    END
  END mem_in_core0[50]
  PIN mem_in_core0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1351.7500 0.5200 1351.8500 ;
    END
  END mem_in_core0[49]
  PIN mem_in_core0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1347.7500 0.5200 1347.8500 ;
    END
  END mem_in_core0[48]
  PIN mem_in_core0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1343.7500 0.5200 1343.8500 ;
    END
  END mem_in_core0[47]
  PIN mem_in_core0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1339.7500 0.5200 1339.8500 ;
    END
  END mem_in_core0[46]
  PIN mem_in_core0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1335.7500 0.5200 1335.8500 ;
    END
  END mem_in_core0[45]
  PIN mem_in_core0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1331.7500 0.5200 1331.8500 ;
    END
  END mem_in_core0[44]
  PIN mem_in_core0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1327.7500 0.5200 1327.8500 ;
    END
  END mem_in_core0[43]
  PIN mem_in_core0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1323.7500 0.5200 1323.8500 ;
    END
  END mem_in_core0[42]
  PIN mem_in_core0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1319.7500 0.5200 1319.8500 ;
    END
  END mem_in_core0[41]
  PIN mem_in_core0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1315.7500 0.5200 1315.8500 ;
    END
  END mem_in_core0[40]
  PIN mem_in_core0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1311.7500 0.5200 1311.8500 ;
    END
  END mem_in_core0[39]
  PIN mem_in_core0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1307.7500 0.5200 1307.8500 ;
    END
  END mem_in_core0[38]
  PIN mem_in_core0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1303.7500 0.5200 1303.8500 ;
    END
  END mem_in_core0[37]
  PIN mem_in_core0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1299.7500 0.5200 1299.8500 ;
    END
  END mem_in_core0[36]
  PIN mem_in_core0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1295.7500 0.5200 1295.8500 ;
    END
  END mem_in_core0[35]
  PIN mem_in_core0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1291.7500 0.5200 1291.8500 ;
    END
  END mem_in_core0[34]
  PIN mem_in_core0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1287.7500 0.5200 1287.8500 ;
    END
  END mem_in_core0[33]
  PIN mem_in_core0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1283.7500 0.5200 1283.8500 ;
    END
  END mem_in_core0[32]
  PIN mem_in_core0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1279.7500 0.5200 1279.8500 ;
    END
  END mem_in_core0[31]
  PIN mem_in_core0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1275.7500 0.5200 1275.8500 ;
    END
  END mem_in_core0[30]
  PIN mem_in_core0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1271.7500 0.5200 1271.8500 ;
    END
  END mem_in_core0[29]
  PIN mem_in_core0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1267.7500 0.5200 1267.8500 ;
    END
  END mem_in_core0[28]
  PIN mem_in_core0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1263.7500 0.5200 1263.8500 ;
    END
  END mem_in_core0[27]
  PIN mem_in_core0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1259.7500 0.5200 1259.8500 ;
    END
  END mem_in_core0[26]
  PIN mem_in_core0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1255.7500 0.5200 1255.8500 ;
    END
  END mem_in_core0[25]
  PIN mem_in_core0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1251.7500 0.5200 1251.8500 ;
    END
  END mem_in_core0[24]
  PIN mem_in_core0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1247.7500 0.5200 1247.8500 ;
    END
  END mem_in_core0[23]
  PIN mem_in_core0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1243.7500 0.5200 1243.8500 ;
    END
  END mem_in_core0[22]
  PIN mem_in_core0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1239.7500 0.5200 1239.8500 ;
    END
  END mem_in_core0[21]
  PIN mem_in_core0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1235.7500 0.5200 1235.8500 ;
    END
  END mem_in_core0[20]
  PIN mem_in_core0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1231.7500 0.5200 1231.8500 ;
    END
  END mem_in_core0[19]
  PIN mem_in_core0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1227.7500 0.5200 1227.8500 ;
    END
  END mem_in_core0[18]
  PIN mem_in_core0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1223.7500 0.5200 1223.8500 ;
    END
  END mem_in_core0[17]
  PIN mem_in_core0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1219.7500 0.5200 1219.8500 ;
    END
  END mem_in_core0[16]
  PIN mem_in_core0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1215.7500 0.5200 1215.8500 ;
    END
  END mem_in_core0[15]
  PIN mem_in_core0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1211.7500 0.5200 1211.8500 ;
    END
  END mem_in_core0[14]
  PIN mem_in_core0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1207.7500 0.5200 1207.8500 ;
    END
  END mem_in_core0[13]
  PIN mem_in_core0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1203.7500 0.5200 1203.8500 ;
    END
  END mem_in_core0[12]
  PIN mem_in_core0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1199.7500 0.5200 1199.8500 ;
    END
  END mem_in_core0[11]
  PIN mem_in_core0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1195.7500 0.5200 1195.8500 ;
    END
  END mem_in_core0[10]
  PIN mem_in_core0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1191.7500 0.5200 1191.8500 ;
    END
  END mem_in_core0[9]
  PIN mem_in_core0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1187.7500 0.5200 1187.8500 ;
    END
  END mem_in_core0[8]
  PIN mem_in_core0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1183.7500 0.5200 1183.8500 ;
    END
  END mem_in_core0[7]
  PIN mem_in_core0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1179.7500 0.5200 1179.8500 ;
    END
  END mem_in_core0[6]
  PIN mem_in_core0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1175.7500 0.5200 1175.8500 ;
    END
  END mem_in_core0[5]
  PIN mem_in_core0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1171.7500 0.5200 1171.8500 ;
    END
  END mem_in_core0[4]
  PIN mem_in_core0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1167.7500 0.5200 1167.8500 ;
    END
  END mem_in_core0[3]
  PIN mem_in_core0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1163.7500 0.5200 1163.8500 ;
    END
  END mem_in_core0[2]
  PIN mem_in_core0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1159.7500 0.5200 1159.8500 ;
    END
  END mem_in_core0[1]
  PIN mem_in_core0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1155.7500 0.5200 1155.8500 ;
    END
  END mem_in_core0[0]
  PIN mem_in_core1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1663.7500 0.5200 1663.8500 ;
    END
  END mem_in_core1[63]
  PIN mem_in_core1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1659.7500 0.5200 1659.8500 ;
    END
  END mem_in_core1[62]
  PIN mem_in_core1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1655.7500 0.5200 1655.8500 ;
    END
  END mem_in_core1[61]
  PIN mem_in_core1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1651.7500 0.5200 1651.8500 ;
    END
  END mem_in_core1[60]
  PIN mem_in_core1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1647.7500 0.5200 1647.8500 ;
    END
  END mem_in_core1[59]
  PIN mem_in_core1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1643.7500 0.5200 1643.8500 ;
    END
  END mem_in_core1[58]
  PIN mem_in_core1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1639.7500 0.5200 1639.8500 ;
    END
  END mem_in_core1[57]
  PIN mem_in_core1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1635.7500 0.5200 1635.8500 ;
    END
  END mem_in_core1[56]
  PIN mem_in_core1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1631.7500 0.5200 1631.8500 ;
    END
  END mem_in_core1[55]
  PIN mem_in_core1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1627.7500 0.5200 1627.8500 ;
    END
  END mem_in_core1[54]
  PIN mem_in_core1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1623.7500 0.5200 1623.8500 ;
    END
  END mem_in_core1[53]
  PIN mem_in_core1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1619.7500 0.5200 1619.8500 ;
    END
  END mem_in_core1[52]
  PIN mem_in_core1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1615.7500 0.5200 1615.8500 ;
    END
  END mem_in_core1[51]
  PIN mem_in_core1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1611.7500 0.5200 1611.8500 ;
    END
  END mem_in_core1[50]
  PIN mem_in_core1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1607.7500 0.5200 1607.8500 ;
    END
  END mem_in_core1[49]
  PIN mem_in_core1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1603.7500 0.5200 1603.8500 ;
    END
  END mem_in_core1[48]
  PIN mem_in_core1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1599.7500 0.5200 1599.8500 ;
    END
  END mem_in_core1[47]
  PIN mem_in_core1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1595.7500 0.5200 1595.8500 ;
    END
  END mem_in_core1[46]
  PIN mem_in_core1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1591.7500 0.5200 1591.8500 ;
    END
  END mem_in_core1[45]
  PIN mem_in_core1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1587.7500 0.5200 1587.8500 ;
    END
  END mem_in_core1[44]
  PIN mem_in_core1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1583.7500 0.5200 1583.8500 ;
    END
  END mem_in_core1[43]
  PIN mem_in_core1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1579.7500 0.5200 1579.8500 ;
    END
  END mem_in_core1[42]
  PIN mem_in_core1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1575.7500 0.5200 1575.8500 ;
    END
  END mem_in_core1[41]
  PIN mem_in_core1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1571.7500 0.5200 1571.8500 ;
    END
  END mem_in_core1[40]
  PIN mem_in_core1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1567.7500 0.5200 1567.8500 ;
    END
  END mem_in_core1[39]
  PIN mem_in_core1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1563.7500 0.5200 1563.8500 ;
    END
  END mem_in_core1[38]
  PIN mem_in_core1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1559.7500 0.5200 1559.8500 ;
    END
  END mem_in_core1[37]
  PIN mem_in_core1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1555.7500 0.5200 1555.8500 ;
    END
  END mem_in_core1[36]
  PIN mem_in_core1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1551.7500 0.5200 1551.8500 ;
    END
  END mem_in_core1[35]
  PIN mem_in_core1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1547.7500 0.5200 1547.8500 ;
    END
  END mem_in_core1[34]
  PIN mem_in_core1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1543.7500 0.5200 1543.8500 ;
    END
  END mem_in_core1[33]
  PIN mem_in_core1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1539.7500 0.5200 1539.8500 ;
    END
  END mem_in_core1[32]
  PIN mem_in_core1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1535.7500 0.5200 1535.8500 ;
    END
  END mem_in_core1[31]
  PIN mem_in_core1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1531.7500 0.5200 1531.8500 ;
    END
  END mem_in_core1[30]
  PIN mem_in_core1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1527.7500 0.5200 1527.8500 ;
    END
  END mem_in_core1[29]
  PIN mem_in_core1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1523.7500 0.5200 1523.8500 ;
    END
  END mem_in_core1[28]
  PIN mem_in_core1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1519.7500 0.5200 1519.8500 ;
    END
  END mem_in_core1[27]
  PIN mem_in_core1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1515.7500 0.5200 1515.8500 ;
    END
  END mem_in_core1[26]
  PIN mem_in_core1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1511.7500 0.5200 1511.8500 ;
    END
  END mem_in_core1[25]
  PIN mem_in_core1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1507.7500 0.5200 1507.8500 ;
    END
  END mem_in_core1[24]
  PIN mem_in_core1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1503.7500 0.5200 1503.8500 ;
    END
  END mem_in_core1[23]
  PIN mem_in_core1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1499.7500 0.5200 1499.8500 ;
    END
  END mem_in_core1[22]
  PIN mem_in_core1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1495.7500 0.5200 1495.8500 ;
    END
  END mem_in_core1[21]
  PIN mem_in_core1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1491.7500 0.5200 1491.8500 ;
    END
  END mem_in_core1[20]
  PIN mem_in_core1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1487.7500 0.5200 1487.8500 ;
    END
  END mem_in_core1[19]
  PIN mem_in_core1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1483.7500 0.5200 1483.8500 ;
    END
  END mem_in_core1[18]
  PIN mem_in_core1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1479.7500 0.5200 1479.8500 ;
    END
  END mem_in_core1[17]
  PIN mem_in_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1475.7500 0.5200 1475.8500 ;
    END
  END mem_in_core1[16]
  PIN mem_in_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1471.7500 0.5200 1471.8500 ;
    END
  END mem_in_core1[15]
  PIN mem_in_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1467.7500 0.5200 1467.8500 ;
    END
  END mem_in_core1[14]
  PIN mem_in_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1463.7500 0.5200 1463.8500 ;
    END
  END mem_in_core1[13]
  PIN mem_in_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1459.7500 0.5200 1459.8500 ;
    END
  END mem_in_core1[12]
  PIN mem_in_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1455.7500 0.5200 1455.8500 ;
    END
  END mem_in_core1[11]
  PIN mem_in_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1451.7500 0.5200 1451.8500 ;
    END
  END mem_in_core1[10]
  PIN mem_in_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1447.7500 0.5200 1447.8500 ;
    END
  END mem_in_core1[9]
  PIN mem_in_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1443.7500 0.5200 1443.8500 ;
    END
  END mem_in_core1[8]
  PIN mem_in_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1439.7500 0.5200 1439.8500 ;
    END
  END mem_in_core1[7]
  PIN mem_in_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1435.7500 0.5200 1435.8500 ;
    END
  END mem_in_core1[6]
  PIN mem_in_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1431.7500 0.5200 1431.8500 ;
    END
  END mem_in_core1[5]
  PIN mem_in_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1427.7500 0.5200 1427.8500 ;
    END
  END mem_in_core1[4]
  PIN mem_in_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1423.7500 0.5200 1423.8500 ;
    END
  END mem_in_core1[3]
  PIN mem_in_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1419.7500 0.5200 1419.8500 ;
    END
  END mem_in_core1[2]
  PIN mem_in_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1415.7500 0.5200 1415.8500 ;
    END
  END mem_in_core1[1]
  PIN mem_in_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1411.7500 0.5200 1411.8500 ;
    END
  END mem_in_core1[0]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1445.7500 0.5200 1445.8500 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1441.7500 0.5200 1441.8500 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1437.7500 0.5200 1437.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1433.7500 0.5200 1433.8500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1429.7500 0.5200 1429.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1425.7500 0.5200 1425.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1421.7500 0.5200 1421.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1417.7500 0.5200 1417.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1413.7500 0.5200 1413.8500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1409.7500 0.5200 1409.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1405.7500 0.5200 1405.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1401.7500 0.5200 1401.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1397.7500 0.5200 1397.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1393.7500 0.5200 1393.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1389.7500 0.5200 1389.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1385.7500 0.5200 1385.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1381.7500 0.5200 1381.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1377.7500 0.5200 1377.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1373.7500 0.5200 1373.8500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1449.7500 0.5200 1449.8500 ;
    END
  END reset
  PIN out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 772.1500 1420.0000 772.2500 ;
    END
  END out[319]
  PIN out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 776.1500 1420.0000 776.2500 ;
    END
  END out[318]
  PIN out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 780.1500 1420.0000 780.2500 ;
    END
  END out[317]
  PIN out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 784.1500 1420.0000 784.2500 ;
    END
  END out[316]
  PIN out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 788.1500 1420.0000 788.2500 ;
    END
  END out[315]
  PIN out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 792.1500 1420.0000 792.2500 ;
    END
  END out[314]
  PIN out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 796.1500 1420.0000 796.2500 ;
    END
  END out[313]
  PIN out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 800.1500 1420.0000 800.2500 ;
    END
  END out[312]
  PIN out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 804.1500 1420.0000 804.2500 ;
    END
  END out[311]
  PIN out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 808.1500 1420.0000 808.2500 ;
    END
  END out[310]
  PIN out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 812.1500 1420.0000 812.2500 ;
    END
  END out[309]
  PIN out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 816.1500 1420.0000 816.2500 ;
    END
  END out[308]
  PIN out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 820.1500 1420.0000 820.2500 ;
    END
  END out[307]
  PIN out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 824.1500 1420.0000 824.2500 ;
    END
  END out[306]
  PIN out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 828.1500 1420.0000 828.2500 ;
    END
  END out[305]
  PIN out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 832.1500 1420.0000 832.2500 ;
    END
  END out[304]
  PIN out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 836.1500 1420.0000 836.2500 ;
    END
  END out[303]
  PIN out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 840.1500 1420.0000 840.2500 ;
    END
  END out[302]
  PIN out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 844.1500 1420.0000 844.2500 ;
    END
  END out[301]
  PIN out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 848.1500 1420.0000 848.2500 ;
    END
  END out[300]
  PIN out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 852.1500 1420.0000 852.2500 ;
    END
  END out[299]
  PIN out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 856.1500 1420.0000 856.2500 ;
    END
  END out[298]
  PIN out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 860.1500 1420.0000 860.2500 ;
    END
  END out[297]
  PIN out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 864.1500 1420.0000 864.2500 ;
    END
  END out[296]
  PIN out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 868.1500 1420.0000 868.2500 ;
    END
  END out[295]
  PIN out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 872.1500 1420.0000 872.2500 ;
    END
  END out[294]
  PIN out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 876.1500 1420.0000 876.2500 ;
    END
  END out[293]
  PIN out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 880.1500 1420.0000 880.2500 ;
    END
  END out[292]
  PIN out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 884.1500 1420.0000 884.2500 ;
    END
  END out[291]
  PIN out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 888.1500 1420.0000 888.2500 ;
    END
  END out[290]
  PIN out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 892.1500 1420.0000 892.2500 ;
    END
  END out[289]
  PIN out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 896.1500 1420.0000 896.2500 ;
    END
  END out[288]
  PIN out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 900.1500 1420.0000 900.2500 ;
    END
  END out[287]
  PIN out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 904.1500 1420.0000 904.2500 ;
    END
  END out[286]
  PIN out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 908.1500 1420.0000 908.2500 ;
    END
  END out[285]
  PIN out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 912.1500 1420.0000 912.2500 ;
    END
  END out[284]
  PIN out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 916.1500 1420.0000 916.2500 ;
    END
  END out[283]
  PIN out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 920.1500 1420.0000 920.2500 ;
    END
  END out[282]
  PIN out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 924.1500 1420.0000 924.2500 ;
    END
  END out[281]
  PIN out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 928.1500 1420.0000 928.2500 ;
    END
  END out[280]
  PIN out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 932.1500 1420.0000 932.2500 ;
    END
  END out[279]
  PIN out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 936.1500 1420.0000 936.2500 ;
    END
  END out[278]
  PIN out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 940.1500 1420.0000 940.2500 ;
    END
  END out[277]
  PIN out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 944.1500 1420.0000 944.2500 ;
    END
  END out[276]
  PIN out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 948.1500 1420.0000 948.2500 ;
    END
  END out[275]
  PIN out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 952.1500 1420.0000 952.2500 ;
    END
  END out[274]
  PIN out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 956.1500 1420.0000 956.2500 ;
    END
  END out[273]
  PIN out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 960.1500 1420.0000 960.2500 ;
    END
  END out[272]
  PIN out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 964.1500 1420.0000 964.2500 ;
    END
  END out[271]
  PIN out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 968.1500 1420.0000 968.2500 ;
    END
  END out[270]
  PIN out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 972.1500 1420.0000 972.2500 ;
    END
  END out[269]
  PIN out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 976.1500 1420.0000 976.2500 ;
    END
  END out[268]
  PIN out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 980.1500 1420.0000 980.2500 ;
    END
  END out[267]
  PIN out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 984.1500 1420.0000 984.2500 ;
    END
  END out[266]
  PIN out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 988.1500 1420.0000 988.2500 ;
    END
  END out[265]
  PIN out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 992.1500 1420.0000 992.2500 ;
    END
  END out[264]
  PIN out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 996.1500 1420.0000 996.2500 ;
    END
  END out[263]
  PIN out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1000.1500 1420.0000 1000.2500 ;
    END
  END out[262]
  PIN out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1004.1500 1420.0000 1004.2500 ;
    END
  END out[261]
  PIN out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1008.1500 1420.0000 1008.2500 ;
    END
  END out[260]
  PIN out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1012.1500 1420.0000 1012.2500 ;
    END
  END out[259]
  PIN out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1016.1500 1420.0000 1016.2500 ;
    END
  END out[258]
  PIN out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1020.1500 1420.0000 1020.2500 ;
    END
  END out[257]
  PIN out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1024.1500 1420.0000 1024.2500 ;
    END
  END out[256]
  PIN out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1028.1500 1420.0000 1028.2500 ;
    END
  END out[255]
  PIN out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1032.1500 1420.0000 1032.2500 ;
    END
  END out[254]
  PIN out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1036.1500 1420.0000 1036.2500 ;
    END
  END out[253]
  PIN out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1040.1500 1420.0000 1040.2500 ;
    END
  END out[252]
  PIN out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1044.1500 1420.0000 1044.2500 ;
    END
  END out[251]
  PIN out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1048.1500 1420.0000 1048.2500 ;
    END
  END out[250]
  PIN out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1052.1500 1420.0000 1052.2500 ;
    END
  END out[249]
  PIN out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1056.1500 1420.0000 1056.2500 ;
    END
  END out[248]
  PIN out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1060.1500 1420.0000 1060.2500 ;
    END
  END out[247]
  PIN out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1064.1500 1420.0000 1064.2500 ;
    END
  END out[246]
  PIN out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1068.1500 1420.0000 1068.2500 ;
    END
  END out[245]
  PIN out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1072.1500 1420.0000 1072.2500 ;
    END
  END out[244]
  PIN out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1076.1500 1420.0000 1076.2500 ;
    END
  END out[243]
  PIN out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1080.1500 1420.0000 1080.2500 ;
    END
  END out[242]
  PIN out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1084.1500 1420.0000 1084.2500 ;
    END
  END out[241]
  PIN out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1088.1500 1420.0000 1088.2500 ;
    END
  END out[240]
  PIN out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1092.1500 1420.0000 1092.2500 ;
    END
  END out[239]
  PIN out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1096.1500 1420.0000 1096.2500 ;
    END
  END out[238]
  PIN out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1100.1500 1420.0000 1100.2500 ;
    END
  END out[237]
  PIN out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1104.1500 1420.0000 1104.2500 ;
    END
  END out[236]
  PIN out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1108.1500 1420.0000 1108.2500 ;
    END
  END out[235]
  PIN out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1112.1500 1420.0000 1112.2500 ;
    END
  END out[234]
  PIN out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1116.1500 1420.0000 1116.2500 ;
    END
  END out[233]
  PIN out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1120.1500 1420.0000 1120.2500 ;
    END
  END out[232]
  PIN out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1124.1500 1420.0000 1124.2500 ;
    END
  END out[231]
  PIN out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1128.1500 1420.0000 1128.2500 ;
    END
  END out[230]
  PIN out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1132.1500 1420.0000 1132.2500 ;
    END
  END out[229]
  PIN out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1136.1500 1420.0000 1136.2500 ;
    END
  END out[228]
  PIN out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1140.1500 1420.0000 1140.2500 ;
    END
  END out[227]
  PIN out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1144.1500 1420.0000 1144.2500 ;
    END
  END out[226]
  PIN out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1148.1500 1420.0000 1148.2500 ;
    END
  END out[225]
  PIN out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1152.1500 1420.0000 1152.2500 ;
    END
  END out[224]
  PIN out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1156.1500 1420.0000 1156.2500 ;
    END
  END out[223]
  PIN out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1160.1500 1420.0000 1160.2500 ;
    END
  END out[222]
  PIN out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1164.1500 1420.0000 1164.2500 ;
    END
  END out[221]
  PIN out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1168.1500 1420.0000 1168.2500 ;
    END
  END out[220]
  PIN out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1172.1500 1420.0000 1172.2500 ;
    END
  END out[219]
  PIN out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1176.1500 1420.0000 1176.2500 ;
    END
  END out[218]
  PIN out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1180.1500 1420.0000 1180.2500 ;
    END
  END out[217]
  PIN out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1184.1500 1420.0000 1184.2500 ;
    END
  END out[216]
  PIN out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1188.1500 1420.0000 1188.2500 ;
    END
  END out[215]
  PIN out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1192.1500 1420.0000 1192.2500 ;
    END
  END out[214]
  PIN out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1196.1500 1420.0000 1196.2500 ;
    END
  END out[213]
  PIN out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1200.1500 1420.0000 1200.2500 ;
    END
  END out[212]
  PIN out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1204.1500 1420.0000 1204.2500 ;
    END
  END out[211]
  PIN out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1208.1500 1420.0000 1208.2500 ;
    END
  END out[210]
  PIN out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1212.1500 1420.0000 1212.2500 ;
    END
  END out[209]
  PIN out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1216.1500 1420.0000 1216.2500 ;
    END
  END out[208]
  PIN out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1220.1500 1420.0000 1220.2500 ;
    END
  END out[207]
  PIN out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1224.1500 1420.0000 1224.2500 ;
    END
  END out[206]
  PIN out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1228.1500 1420.0000 1228.2500 ;
    END
  END out[205]
  PIN out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1232.1500 1420.0000 1232.2500 ;
    END
  END out[204]
  PIN out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1236.1500 1420.0000 1236.2500 ;
    END
  END out[203]
  PIN out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1240.1500 1420.0000 1240.2500 ;
    END
  END out[202]
  PIN out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1244.1500 1420.0000 1244.2500 ;
    END
  END out[201]
  PIN out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1248.1500 1420.0000 1248.2500 ;
    END
  END out[200]
  PIN out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1252.1500 1420.0000 1252.2500 ;
    END
  END out[199]
  PIN out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1256.1500 1420.0000 1256.2500 ;
    END
  END out[198]
  PIN out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1260.1500 1420.0000 1260.2500 ;
    END
  END out[197]
  PIN out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1264.1500 1420.0000 1264.2500 ;
    END
  END out[196]
  PIN out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1268.1500 1420.0000 1268.2500 ;
    END
  END out[195]
  PIN out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1272.1500 1420.0000 1272.2500 ;
    END
  END out[194]
  PIN out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1276.1500 1420.0000 1276.2500 ;
    END
  END out[193]
  PIN out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1280.1500 1420.0000 1280.2500 ;
    END
  END out[192]
  PIN out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1284.1500 1420.0000 1284.2500 ;
    END
  END out[191]
  PIN out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1288.1500 1420.0000 1288.2500 ;
    END
  END out[190]
  PIN out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1292.1500 1420.0000 1292.2500 ;
    END
  END out[189]
  PIN out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1296.1500 1420.0000 1296.2500 ;
    END
  END out[188]
  PIN out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1300.1500 1420.0000 1300.2500 ;
    END
  END out[187]
  PIN out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1304.1500 1420.0000 1304.2500 ;
    END
  END out[186]
  PIN out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1308.1500 1420.0000 1308.2500 ;
    END
  END out[185]
  PIN out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1312.1500 1420.0000 1312.2500 ;
    END
  END out[184]
  PIN out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1316.1500 1420.0000 1316.2500 ;
    END
  END out[183]
  PIN out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1320.1500 1420.0000 1320.2500 ;
    END
  END out[182]
  PIN out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1324.1500 1420.0000 1324.2500 ;
    END
  END out[181]
  PIN out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1328.1500 1420.0000 1328.2500 ;
    END
  END out[180]
  PIN out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1332.1500 1420.0000 1332.2500 ;
    END
  END out[179]
  PIN out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1336.1500 1420.0000 1336.2500 ;
    END
  END out[178]
  PIN out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1340.1500 1420.0000 1340.2500 ;
    END
  END out[177]
  PIN out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1344.1500 1420.0000 1344.2500 ;
    END
  END out[176]
  PIN out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1348.1500 1420.0000 1348.2500 ;
    END
  END out[175]
  PIN out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1352.1500 1420.0000 1352.2500 ;
    END
  END out[174]
  PIN out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1356.1500 1420.0000 1356.2500 ;
    END
  END out[173]
  PIN out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1360.1500 1420.0000 1360.2500 ;
    END
  END out[172]
  PIN out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1364.1500 1420.0000 1364.2500 ;
    END
  END out[171]
  PIN out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1368.1500 1420.0000 1368.2500 ;
    END
  END out[170]
  PIN out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1372.1500 1420.0000 1372.2500 ;
    END
  END out[169]
  PIN out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1376.1500 1420.0000 1376.2500 ;
    END
  END out[168]
  PIN out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1380.1500 1420.0000 1380.2500 ;
    END
  END out[167]
  PIN out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1384.1500 1420.0000 1384.2500 ;
    END
  END out[166]
  PIN out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1388.1500 1420.0000 1388.2500 ;
    END
  END out[165]
  PIN out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1392.1500 1420.0000 1392.2500 ;
    END
  END out[164]
  PIN out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1396.1500 1420.0000 1396.2500 ;
    END
  END out[163]
  PIN out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1400.1500 1420.0000 1400.2500 ;
    END
  END out[162]
  PIN out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1404.1500 1420.0000 1404.2500 ;
    END
  END out[161]
  PIN out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1408.1500 1420.0000 1408.2500 ;
    END
  END out[160]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1412.1500 1420.0000 1412.2500 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1416.1500 1420.0000 1416.2500 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1420.1500 1420.0000 1420.2500 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1424.1500 1420.0000 1424.2500 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1428.1500 1420.0000 1428.2500 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1432.1500 1420.0000 1432.2500 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1436.1500 1420.0000 1436.2500 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1440.1500 1420.0000 1440.2500 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1444.1500 1420.0000 1444.2500 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1448.1500 1420.0000 1448.2500 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1452.1500 1420.0000 1452.2500 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1456.1500 1420.0000 1456.2500 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1460.1500 1420.0000 1460.2500 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1464.1500 1420.0000 1464.2500 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1468.1500 1420.0000 1468.2500 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1472.1500 1420.0000 1472.2500 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1476.1500 1420.0000 1476.2500 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1480.1500 1420.0000 1480.2500 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1484.1500 1420.0000 1484.2500 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1488.1500 1420.0000 1488.2500 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1492.1500 1420.0000 1492.2500 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1496.1500 1420.0000 1496.2500 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1500.1500 1420.0000 1500.2500 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1504.1500 1420.0000 1504.2500 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1508.1500 1420.0000 1508.2500 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1512.1500 1420.0000 1512.2500 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1516.1500 1420.0000 1516.2500 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1520.1500 1420.0000 1520.2500 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1524.1500 1420.0000 1524.2500 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1528.1500 1420.0000 1528.2500 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1532.1500 1420.0000 1532.2500 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1536.1500 1420.0000 1536.2500 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1540.1500 1420.0000 1540.2500 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1544.1500 1420.0000 1544.2500 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1548.1500 1420.0000 1548.2500 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1552.1500 1420.0000 1552.2500 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1556.1500 1420.0000 1556.2500 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1560.1500 1420.0000 1560.2500 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1564.1500 1420.0000 1564.2500 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1568.1500 1420.0000 1568.2500 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1572.1500 1420.0000 1572.2500 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1576.1500 1420.0000 1576.2500 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1580.1500 1420.0000 1580.2500 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1584.1500 1420.0000 1584.2500 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1588.1500 1420.0000 1588.2500 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1592.1500 1420.0000 1592.2500 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1596.1500 1420.0000 1596.2500 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1600.1500 1420.0000 1600.2500 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1604.1500 1420.0000 1604.2500 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1608.1500 1420.0000 1608.2500 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1612.1500 1420.0000 1612.2500 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1616.1500 1420.0000 1616.2500 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1620.1500 1420.0000 1620.2500 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1624.1500 1420.0000 1624.2500 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1628.1500 1420.0000 1628.2500 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1632.1500 1420.0000 1632.2500 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1636.1500 1420.0000 1636.2500 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1640.1500 1420.0000 1640.2500 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1644.1500 1420.0000 1644.2500 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1648.1500 1420.0000 1648.2500 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1652.1500 1420.0000 1652.2500 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1656.1500 1420.0000 1656.2500 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1660.1500 1420.0000 1660.2500 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1664.1500 1420.0000 1664.2500 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1668.1500 1420.0000 1668.2500 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1672.1500 1420.0000 1672.2500 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1676.1500 1420.0000 1676.2500 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1680.1500 1420.0000 1680.2500 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1684.1500 1420.0000 1684.2500 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1688.1500 1420.0000 1688.2500 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1692.1500 1420.0000 1692.2500 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1696.1500 1420.0000 1696.2500 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1700.1500 1420.0000 1700.2500 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1704.1500 1420.0000 1704.2500 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1708.1500 1420.0000 1708.2500 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1712.1500 1420.0000 1712.2500 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1716.1500 1420.0000 1716.2500 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1720.1500 1420.0000 1720.2500 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1724.1500 1420.0000 1724.2500 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1728.1500 1420.0000 1728.2500 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1732.1500 1420.0000 1732.2500 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1736.1500 1420.0000 1736.2500 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1740.1500 1420.0000 1740.2500 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1744.1500 1420.0000 1744.2500 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1748.1500 1420.0000 1748.2500 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1752.1500 1420.0000 1752.2500 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1756.1500 1420.0000 1756.2500 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1760.1500 1420.0000 1760.2500 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1764.1500 1420.0000 1764.2500 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1768.1500 1420.0000 1768.2500 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1772.1500 1420.0000 1772.2500 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1776.1500 1420.0000 1776.2500 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1780.1500 1420.0000 1780.2500 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1784.1500 1420.0000 1784.2500 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1788.1500 1420.0000 1788.2500 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1792.1500 1420.0000 1792.2500 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1796.1500 1420.0000 1796.2500 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1800.1500 1420.0000 1800.2500 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1804.1500 1420.0000 1804.2500 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1808.1500 1420.0000 1808.2500 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1812.1500 1420.0000 1812.2500 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1816.1500 1420.0000 1816.2500 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1820.1500 1420.0000 1820.2500 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1824.1500 1420.0000 1824.2500 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1828.1500 1420.0000 1828.2500 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1832.1500 1420.0000 1832.2500 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1836.1500 1420.0000 1836.2500 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1840.1500 1420.0000 1840.2500 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1844.1500 1420.0000 1844.2500 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1848.1500 1420.0000 1848.2500 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1852.1500 1420.0000 1852.2500 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1856.1500 1420.0000 1856.2500 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1860.1500 1420.0000 1860.2500 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1864.1500 1420.0000 1864.2500 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1868.1500 1420.0000 1868.2500 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1872.1500 1420.0000 1872.2500 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1876.1500 1420.0000 1876.2500 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1880.1500 1420.0000 1880.2500 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1884.1500 1420.0000 1884.2500 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1888.1500 1420.0000 1888.2500 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1892.1500 1420.0000 1892.2500 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1896.1500 1420.0000 1896.2500 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1900.1500 1420.0000 1900.2500 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1904.1500 1420.0000 1904.2500 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1908.1500 1420.0000 1908.2500 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1912.1500 1420.0000 1912.2500 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1916.1500 1420.0000 1916.2500 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1920.1500 1420.0000 1920.2500 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1924.1500 1420.0000 1924.2500 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1928.1500 1420.0000 1928.2500 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1932.1500 1420.0000 1932.2500 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1936.1500 1420.0000 1936.2500 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1940.1500 1420.0000 1940.2500 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1944.1500 1420.0000 1944.2500 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1948.1500 1420.0000 1948.2500 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1952.1500 1420.0000 1952.2500 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1956.1500 1420.0000 1956.2500 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1960.1500 1420.0000 1960.2500 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1964.1500 1420.0000 1964.2500 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1968.1500 1420.0000 1968.2500 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1972.1500 1420.0000 1972.2500 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1976.1500 1420.0000 1976.2500 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1980.1500 1420.0000 1980.2500 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1984.1500 1420.0000 1984.2500 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1988.1500 1420.0000 1988.2500 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1992.1500 1420.0000 1992.2500 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 1996.1500 1420.0000 1996.2500 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2000.1500 1420.0000 2000.2500 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2004.1500 1420.0000 2004.2500 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2008.1500 1420.0000 2008.2500 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2012.1500 1420.0000 2012.2500 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2016.1500 1420.0000 2016.2500 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2020.1500 1420.0000 2020.2500 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2024.1500 1420.0000 2024.2500 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2028.1500 1420.0000 2028.2500 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2032.1500 1420.0000 2032.2500 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2036.1500 1420.0000 2036.2500 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2040.1500 1420.0000 2040.2500 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2044.1500 1420.0000 2044.2500 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1419.4800 2048.1500 1420.0000 2048.2500 ;
    END
  END out[0]
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M3 ;
      RECT 0.0000 2048.3500 1420.0000 2820.0000 ;
      RECT 0.0000 2048.0500 1419.3800 2048.3500 ;
      RECT 0.0000 2044.3500 1420.0000 2048.0500 ;
      RECT 0.0000 2044.0500 1419.3800 2044.3500 ;
      RECT 0.0000 2040.3500 1420.0000 2044.0500 ;
      RECT 0.0000 2040.0500 1419.3800 2040.3500 ;
      RECT 0.0000 2036.3500 1420.0000 2040.0500 ;
      RECT 0.0000 2036.0500 1419.3800 2036.3500 ;
      RECT 0.0000 2032.3500 1420.0000 2036.0500 ;
      RECT 0.0000 2032.0500 1419.3800 2032.3500 ;
      RECT 0.0000 2028.3500 1420.0000 2032.0500 ;
      RECT 0.0000 2028.0500 1419.3800 2028.3500 ;
      RECT 0.0000 2024.3500 1420.0000 2028.0500 ;
      RECT 0.0000 2024.0500 1419.3800 2024.3500 ;
      RECT 0.0000 2020.3500 1420.0000 2024.0500 ;
      RECT 0.0000 2020.0500 1419.3800 2020.3500 ;
      RECT 0.0000 2016.3500 1420.0000 2020.0500 ;
      RECT 0.0000 2016.0500 1419.3800 2016.3500 ;
      RECT 0.0000 2012.3500 1420.0000 2016.0500 ;
      RECT 0.0000 2012.0500 1419.3800 2012.3500 ;
      RECT 0.0000 2008.3500 1420.0000 2012.0500 ;
      RECT 0.0000 2008.0500 1419.3800 2008.3500 ;
      RECT 0.0000 2004.3500 1420.0000 2008.0500 ;
      RECT 0.0000 2004.0500 1419.3800 2004.3500 ;
      RECT 0.0000 2000.3500 1420.0000 2004.0500 ;
      RECT 0.0000 2000.0500 1419.3800 2000.3500 ;
      RECT 0.0000 1996.3500 1420.0000 2000.0500 ;
      RECT 0.0000 1996.0500 1419.3800 1996.3500 ;
      RECT 0.0000 1992.3500 1420.0000 1996.0500 ;
      RECT 0.0000 1992.0500 1419.3800 1992.3500 ;
      RECT 0.0000 1988.3500 1420.0000 1992.0500 ;
      RECT 0.0000 1988.0500 1419.3800 1988.3500 ;
      RECT 0.0000 1984.3500 1420.0000 1988.0500 ;
      RECT 0.0000 1984.0500 1419.3800 1984.3500 ;
      RECT 0.0000 1980.3500 1420.0000 1984.0500 ;
      RECT 0.0000 1980.0500 1419.3800 1980.3500 ;
      RECT 0.0000 1976.3500 1420.0000 1980.0500 ;
      RECT 0.0000 1976.0500 1419.3800 1976.3500 ;
      RECT 0.0000 1972.3500 1420.0000 1976.0500 ;
      RECT 0.0000 1972.0500 1419.3800 1972.3500 ;
      RECT 0.0000 1968.3500 1420.0000 1972.0500 ;
      RECT 0.0000 1968.0500 1419.3800 1968.3500 ;
      RECT 0.0000 1964.3500 1420.0000 1968.0500 ;
      RECT 0.0000 1964.0500 1419.3800 1964.3500 ;
      RECT 0.0000 1960.3500 1420.0000 1964.0500 ;
      RECT 0.0000 1960.0500 1419.3800 1960.3500 ;
      RECT 0.0000 1956.3500 1420.0000 1960.0500 ;
      RECT 0.0000 1956.0500 1419.3800 1956.3500 ;
      RECT 0.0000 1952.3500 1420.0000 1956.0500 ;
      RECT 0.0000 1952.0500 1419.3800 1952.3500 ;
      RECT 0.0000 1948.3500 1420.0000 1952.0500 ;
      RECT 0.0000 1948.0500 1419.3800 1948.3500 ;
      RECT 0.0000 1944.3500 1420.0000 1948.0500 ;
      RECT 0.0000 1944.0500 1419.3800 1944.3500 ;
      RECT 0.0000 1940.3500 1420.0000 1944.0500 ;
      RECT 0.0000 1940.0500 1419.3800 1940.3500 ;
      RECT 0.0000 1936.3500 1420.0000 1940.0500 ;
      RECT 0.0000 1936.0500 1419.3800 1936.3500 ;
      RECT 0.0000 1932.3500 1420.0000 1936.0500 ;
      RECT 0.0000 1932.0500 1419.3800 1932.3500 ;
      RECT 0.0000 1928.3500 1420.0000 1932.0500 ;
      RECT 0.0000 1928.0500 1419.3800 1928.3500 ;
      RECT 0.0000 1924.3500 1420.0000 1928.0500 ;
      RECT 0.0000 1924.0500 1419.3800 1924.3500 ;
      RECT 0.0000 1920.3500 1420.0000 1924.0500 ;
      RECT 0.0000 1920.0500 1419.3800 1920.3500 ;
      RECT 0.0000 1916.3500 1420.0000 1920.0500 ;
      RECT 0.0000 1916.0500 1419.3800 1916.3500 ;
      RECT 0.0000 1912.3500 1420.0000 1916.0500 ;
      RECT 0.0000 1912.0500 1419.3800 1912.3500 ;
      RECT 0.0000 1908.3500 1420.0000 1912.0500 ;
      RECT 0.0000 1908.0500 1419.3800 1908.3500 ;
      RECT 0.0000 1904.3500 1420.0000 1908.0500 ;
      RECT 0.0000 1904.0500 1419.3800 1904.3500 ;
      RECT 0.0000 1900.3500 1420.0000 1904.0500 ;
      RECT 0.0000 1900.0500 1419.3800 1900.3500 ;
      RECT 0.0000 1896.3500 1420.0000 1900.0500 ;
      RECT 0.0000 1896.0500 1419.3800 1896.3500 ;
      RECT 0.0000 1892.3500 1420.0000 1896.0500 ;
      RECT 0.0000 1892.0500 1419.3800 1892.3500 ;
      RECT 0.0000 1888.3500 1420.0000 1892.0500 ;
      RECT 0.0000 1888.0500 1419.3800 1888.3500 ;
      RECT 0.0000 1884.3500 1420.0000 1888.0500 ;
      RECT 0.0000 1884.0500 1419.3800 1884.3500 ;
      RECT 0.0000 1880.3500 1420.0000 1884.0500 ;
      RECT 0.0000 1880.0500 1419.3800 1880.3500 ;
      RECT 0.0000 1876.3500 1420.0000 1880.0500 ;
      RECT 0.0000 1876.0500 1419.3800 1876.3500 ;
      RECT 0.0000 1872.3500 1420.0000 1876.0500 ;
      RECT 0.0000 1872.0500 1419.3800 1872.3500 ;
      RECT 0.0000 1868.3500 1420.0000 1872.0500 ;
      RECT 0.0000 1868.0500 1419.3800 1868.3500 ;
      RECT 0.0000 1864.3500 1420.0000 1868.0500 ;
      RECT 0.0000 1864.0500 1419.3800 1864.3500 ;
      RECT 0.0000 1860.3500 1420.0000 1864.0500 ;
      RECT 0.0000 1860.0500 1419.3800 1860.3500 ;
      RECT 0.0000 1856.3500 1420.0000 1860.0500 ;
      RECT 0.0000 1856.0500 1419.3800 1856.3500 ;
      RECT 0.0000 1852.3500 1420.0000 1856.0500 ;
      RECT 0.0000 1852.0500 1419.3800 1852.3500 ;
      RECT 0.0000 1848.3500 1420.0000 1852.0500 ;
      RECT 0.0000 1848.0500 1419.3800 1848.3500 ;
      RECT 0.0000 1844.3500 1420.0000 1848.0500 ;
      RECT 0.0000 1844.0500 1419.3800 1844.3500 ;
      RECT 0.0000 1840.3500 1420.0000 1844.0500 ;
      RECT 0.0000 1840.0500 1419.3800 1840.3500 ;
      RECT 0.0000 1836.3500 1420.0000 1840.0500 ;
      RECT 0.0000 1836.0500 1419.3800 1836.3500 ;
      RECT 0.0000 1832.3500 1420.0000 1836.0500 ;
      RECT 0.0000 1832.0500 1419.3800 1832.3500 ;
      RECT 0.0000 1828.3500 1420.0000 1832.0500 ;
      RECT 0.0000 1828.0500 1419.3800 1828.3500 ;
      RECT 0.0000 1824.3500 1420.0000 1828.0500 ;
      RECT 0.0000 1824.0500 1419.3800 1824.3500 ;
      RECT 0.0000 1820.3500 1420.0000 1824.0500 ;
      RECT 0.0000 1820.0500 1419.3800 1820.3500 ;
      RECT 0.0000 1816.3500 1420.0000 1820.0500 ;
      RECT 0.0000 1816.0500 1419.3800 1816.3500 ;
      RECT 0.0000 1812.3500 1420.0000 1816.0500 ;
      RECT 0.0000 1812.0500 1419.3800 1812.3500 ;
      RECT 0.0000 1808.3500 1420.0000 1812.0500 ;
      RECT 0.0000 1808.0500 1419.3800 1808.3500 ;
      RECT 0.0000 1804.3500 1420.0000 1808.0500 ;
      RECT 0.0000 1804.0500 1419.3800 1804.3500 ;
      RECT 0.0000 1800.3500 1420.0000 1804.0500 ;
      RECT 0.0000 1800.0500 1419.3800 1800.3500 ;
      RECT 0.0000 1796.3500 1420.0000 1800.0500 ;
      RECT 0.0000 1796.0500 1419.3800 1796.3500 ;
      RECT 0.0000 1792.3500 1420.0000 1796.0500 ;
      RECT 0.0000 1792.0500 1419.3800 1792.3500 ;
      RECT 0.0000 1788.3500 1420.0000 1792.0500 ;
      RECT 0.0000 1788.0500 1419.3800 1788.3500 ;
      RECT 0.0000 1784.3500 1420.0000 1788.0500 ;
      RECT 0.0000 1784.0500 1419.3800 1784.3500 ;
      RECT 0.0000 1780.3500 1420.0000 1784.0500 ;
      RECT 0.0000 1780.0500 1419.3800 1780.3500 ;
      RECT 0.0000 1776.3500 1420.0000 1780.0500 ;
      RECT 0.0000 1776.0500 1419.3800 1776.3500 ;
      RECT 0.0000 1772.3500 1420.0000 1776.0500 ;
      RECT 0.0000 1772.0500 1419.3800 1772.3500 ;
      RECT 0.0000 1768.3500 1420.0000 1772.0500 ;
      RECT 0.0000 1768.0500 1419.3800 1768.3500 ;
      RECT 0.0000 1764.3500 1420.0000 1768.0500 ;
      RECT 0.0000 1764.0500 1419.3800 1764.3500 ;
      RECT 0.0000 1760.3500 1420.0000 1764.0500 ;
      RECT 0.0000 1760.0500 1419.3800 1760.3500 ;
      RECT 0.0000 1756.3500 1420.0000 1760.0500 ;
      RECT 0.0000 1756.0500 1419.3800 1756.3500 ;
      RECT 0.0000 1752.3500 1420.0000 1756.0500 ;
      RECT 0.0000 1752.0500 1419.3800 1752.3500 ;
      RECT 0.0000 1748.3500 1420.0000 1752.0500 ;
      RECT 0.0000 1748.0500 1419.3800 1748.3500 ;
      RECT 0.0000 1744.3500 1420.0000 1748.0500 ;
      RECT 0.0000 1744.0500 1419.3800 1744.3500 ;
      RECT 0.0000 1740.3500 1420.0000 1744.0500 ;
      RECT 0.0000 1740.0500 1419.3800 1740.3500 ;
      RECT 0.0000 1736.3500 1420.0000 1740.0500 ;
      RECT 0.0000 1736.0500 1419.3800 1736.3500 ;
      RECT 0.0000 1732.3500 1420.0000 1736.0500 ;
      RECT 0.0000 1732.0500 1419.3800 1732.3500 ;
      RECT 0.0000 1728.3500 1420.0000 1732.0500 ;
      RECT 0.0000 1728.0500 1419.3800 1728.3500 ;
      RECT 0.0000 1724.3500 1420.0000 1728.0500 ;
      RECT 0.0000 1724.0500 1419.3800 1724.3500 ;
      RECT 0.0000 1720.3500 1420.0000 1724.0500 ;
      RECT 0.0000 1720.0500 1419.3800 1720.3500 ;
      RECT 0.0000 1716.3500 1420.0000 1720.0500 ;
      RECT 0.0000 1716.0500 1419.3800 1716.3500 ;
      RECT 0.0000 1712.3500 1420.0000 1716.0500 ;
      RECT 0.0000 1712.0500 1419.3800 1712.3500 ;
      RECT 0.0000 1708.3500 1420.0000 1712.0500 ;
      RECT 0.0000 1708.0500 1419.3800 1708.3500 ;
      RECT 0.0000 1704.3500 1420.0000 1708.0500 ;
      RECT 0.0000 1704.0500 1419.3800 1704.3500 ;
      RECT 0.0000 1700.3500 1420.0000 1704.0500 ;
      RECT 0.0000 1700.0500 1419.3800 1700.3500 ;
      RECT 0.0000 1696.3500 1420.0000 1700.0500 ;
      RECT 0.0000 1696.0500 1419.3800 1696.3500 ;
      RECT 0.0000 1692.3500 1420.0000 1696.0500 ;
      RECT 0.0000 1692.0500 1419.3800 1692.3500 ;
      RECT 0.0000 1688.3500 1420.0000 1692.0500 ;
      RECT 0.0000 1688.0500 1419.3800 1688.3500 ;
      RECT 0.0000 1684.3500 1420.0000 1688.0500 ;
      RECT 0.0000 1684.0500 1419.3800 1684.3500 ;
      RECT 0.0000 1680.3500 1420.0000 1684.0500 ;
      RECT 0.0000 1680.0500 1419.3800 1680.3500 ;
      RECT 0.0000 1676.3500 1420.0000 1680.0500 ;
      RECT 0.0000 1676.0500 1419.3800 1676.3500 ;
      RECT 0.0000 1672.3500 1420.0000 1676.0500 ;
      RECT 0.0000 1672.0500 1419.3800 1672.3500 ;
      RECT 0.0000 1668.3500 1420.0000 1672.0500 ;
      RECT 0.0000 1668.0500 1419.3800 1668.3500 ;
      RECT 0.0000 1664.3500 1420.0000 1668.0500 ;
      RECT 0.0000 1664.0500 1419.3800 1664.3500 ;
      RECT 0.0000 1663.9500 1420.0000 1664.0500 ;
      RECT 0.6200 1663.6500 1420.0000 1663.9500 ;
      RECT 0.0000 1660.3500 1420.0000 1663.6500 ;
      RECT 0.0000 1660.0500 1419.3800 1660.3500 ;
      RECT 0.0000 1659.9500 1420.0000 1660.0500 ;
      RECT 0.6200 1659.6500 1420.0000 1659.9500 ;
      RECT 0.0000 1656.3500 1420.0000 1659.6500 ;
      RECT 0.0000 1656.0500 1419.3800 1656.3500 ;
      RECT 0.0000 1655.9500 1420.0000 1656.0500 ;
      RECT 0.6200 1655.6500 1420.0000 1655.9500 ;
      RECT 0.0000 1652.3500 1420.0000 1655.6500 ;
      RECT 0.0000 1652.0500 1419.3800 1652.3500 ;
      RECT 0.0000 1651.9500 1420.0000 1652.0500 ;
      RECT 0.6200 1651.6500 1420.0000 1651.9500 ;
      RECT 0.0000 1648.3500 1420.0000 1651.6500 ;
      RECT 0.0000 1648.0500 1419.3800 1648.3500 ;
      RECT 0.0000 1647.9500 1420.0000 1648.0500 ;
      RECT 0.6200 1647.6500 1420.0000 1647.9500 ;
      RECT 0.0000 1644.3500 1420.0000 1647.6500 ;
      RECT 0.0000 1644.0500 1419.3800 1644.3500 ;
      RECT 0.0000 1643.9500 1420.0000 1644.0500 ;
      RECT 0.6200 1643.6500 1420.0000 1643.9500 ;
      RECT 0.0000 1640.3500 1420.0000 1643.6500 ;
      RECT 0.0000 1640.0500 1419.3800 1640.3500 ;
      RECT 0.0000 1639.9500 1420.0000 1640.0500 ;
      RECT 0.6200 1639.6500 1420.0000 1639.9500 ;
      RECT 0.0000 1636.3500 1420.0000 1639.6500 ;
      RECT 0.0000 1636.0500 1419.3800 1636.3500 ;
      RECT 0.0000 1635.9500 1420.0000 1636.0500 ;
      RECT 0.6200 1635.6500 1420.0000 1635.9500 ;
      RECT 0.0000 1632.3500 1420.0000 1635.6500 ;
      RECT 0.0000 1632.0500 1419.3800 1632.3500 ;
      RECT 0.0000 1631.9500 1420.0000 1632.0500 ;
      RECT 0.6200 1631.6500 1420.0000 1631.9500 ;
      RECT 0.0000 1628.3500 1420.0000 1631.6500 ;
      RECT 0.0000 1628.0500 1419.3800 1628.3500 ;
      RECT 0.0000 1627.9500 1420.0000 1628.0500 ;
      RECT 0.6200 1627.6500 1420.0000 1627.9500 ;
      RECT 0.0000 1624.3500 1420.0000 1627.6500 ;
      RECT 0.0000 1624.0500 1419.3800 1624.3500 ;
      RECT 0.0000 1623.9500 1420.0000 1624.0500 ;
      RECT 0.6200 1623.6500 1420.0000 1623.9500 ;
      RECT 0.0000 1620.3500 1420.0000 1623.6500 ;
      RECT 0.0000 1620.0500 1419.3800 1620.3500 ;
      RECT 0.0000 1619.9500 1420.0000 1620.0500 ;
      RECT 0.6200 1619.6500 1420.0000 1619.9500 ;
      RECT 0.0000 1616.3500 1420.0000 1619.6500 ;
      RECT 0.0000 1616.0500 1419.3800 1616.3500 ;
      RECT 0.0000 1615.9500 1420.0000 1616.0500 ;
      RECT 0.6200 1615.6500 1420.0000 1615.9500 ;
      RECT 0.0000 1612.3500 1420.0000 1615.6500 ;
      RECT 0.0000 1612.0500 1419.3800 1612.3500 ;
      RECT 0.0000 1611.9500 1420.0000 1612.0500 ;
      RECT 0.6200 1611.6500 1420.0000 1611.9500 ;
      RECT 0.0000 1608.3500 1420.0000 1611.6500 ;
      RECT 0.0000 1608.0500 1419.3800 1608.3500 ;
      RECT 0.0000 1607.9500 1420.0000 1608.0500 ;
      RECT 0.6200 1607.6500 1420.0000 1607.9500 ;
      RECT 0.0000 1604.3500 1420.0000 1607.6500 ;
      RECT 0.0000 1604.0500 1419.3800 1604.3500 ;
      RECT 0.0000 1603.9500 1420.0000 1604.0500 ;
      RECT 0.6200 1603.6500 1420.0000 1603.9500 ;
      RECT 0.0000 1600.3500 1420.0000 1603.6500 ;
      RECT 0.0000 1600.0500 1419.3800 1600.3500 ;
      RECT 0.0000 1599.9500 1420.0000 1600.0500 ;
      RECT 0.6200 1599.6500 1420.0000 1599.9500 ;
      RECT 0.0000 1596.3500 1420.0000 1599.6500 ;
      RECT 0.0000 1596.0500 1419.3800 1596.3500 ;
      RECT 0.0000 1595.9500 1420.0000 1596.0500 ;
      RECT 0.6200 1595.6500 1420.0000 1595.9500 ;
      RECT 0.0000 1592.3500 1420.0000 1595.6500 ;
      RECT 0.0000 1592.0500 1419.3800 1592.3500 ;
      RECT 0.0000 1591.9500 1420.0000 1592.0500 ;
      RECT 0.6200 1591.6500 1420.0000 1591.9500 ;
      RECT 0.0000 1588.3500 1420.0000 1591.6500 ;
      RECT 0.0000 1588.0500 1419.3800 1588.3500 ;
      RECT 0.0000 1587.9500 1420.0000 1588.0500 ;
      RECT 0.6200 1587.6500 1420.0000 1587.9500 ;
      RECT 0.0000 1584.3500 1420.0000 1587.6500 ;
      RECT 0.0000 1584.0500 1419.3800 1584.3500 ;
      RECT 0.0000 1583.9500 1420.0000 1584.0500 ;
      RECT 0.6200 1583.6500 1420.0000 1583.9500 ;
      RECT 0.0000 1580.3500 1420.0000 1583.6500 ;
      RECT 0.0000 1580.0500 1419.3800 1580.3500 ;
      RECT 0.0000 1579.9500 1420.0000 1580.0500 ;
      RECT 0.6200 1579.6500 1420.0000 1579.9500 ;
      RECT 0.0000 1576.3500 1420.0000 1579.6500 ;
      RECT 0.0000 1576.0500 1419.3800 1576.3500 ;
      RECT 0.0000 1575.9500 1420.0000 1576.0500 ;
      RECT 0.6200 1575.6500 1420.0000 1575.9500 ;
      RECT 0.0000 1572.3500 1420.0000 1575.6500 ;
      RECT 0.0000 1572.0500 1419.3800 1572.3500 ;
      RECT 0.0000 1571.9500 1420.0000 1572.0500 ;
      RECT 0.6200 1571.6500 1420.0000 1571.9500 ;
      RECT 0.0000 1568.3500 1420.0000 1571.6500 ;
      RECT 0.0000 1568.0500 1419.3800 1568.3500 ;
      RECT 0.0000 1567.9500 1420.0000 1568.0500 ;
      RECT 0.6200 1567.6500 1420.0000 1567.9500 ;
      RECT 0.0000 1564.3500 1420.0000 1567.6500 ;
      RECT 0.0000 1564.0500 1419.3800 1564.3500 ;
      RECT 0.0000 1563.9500 1420.0000 1564.0500 ;
      RECT 0.6200 1563.6500 1420.0000 1563.9500 ;
      RECT 0.0000 1560.3500 1420.0000 1563.6500 ;
      RECT 0.0000 1560.0500 1419.3800 1560.3500 ;
      RECT 0.0000 1559.9500 1420.0000 1560.0500 ;
      RECT 0.6200 1559.6500 1420.0000 1559.9500 ;
      RECT 0.0000 1556.3500 1420.0000 1559.6500 ;
      RECT 0.0000 1556.0500 1419.3800 1556.3500 ;
      RECT 0.0000 1555.9500 1420.0000 1556.0500 ;
      RECT 0.6200 1555.6500 1420.0000 1555.9500 ;
      RECT 0.0000 1552.3500 1420.0000 1555.6500 ;
      RECT 0.0000 1552.0500 1419.3800 1552.3500 ;
      RECT 0.0000 1551.9500 1420.0000 1552.0500 ;
      RECT 0.6200 1551.6500 1420.0000 1551.9500 ;
      RECT 0.0000 1548.3500 1420.0000 1551.6500 ;
      RECT 0.0000 1548.0500 1419.3800 1548.3500 ;
      RECT 0.0000 1547.9500 1420.0000 1548.0500 ;
      RECT 0.6200 1547.6500 1420.0000 1547.9500 ;
      RECT 0.0000 1544.3500 1420.0000 1547.6500 ;
      RECT 0.0000 1544.0500 1419.3800 1544.3500 ;
      RECT 0.0000 1543.9500 1420.0000 1544.0500 ;
      RECT 0.6200 1543.6500 1420.0000 1543.9500 ;
      RECT 0.0000 1540.3500 1420.0000 1543.6500 ;
      RECT 0.0000 1540.0500 1419.3800 1540.3500 ;
      RECT 0.0000 1539.9500 1420.0000 1540.0500 ;
      RECT 0.6200 1539.6500 1420.0000 1539.9500 ;
      RECT 0.0000 1536.3500 1420.0000 1539.6500 ;
      RECT 0.0000 1536.0500 1419.3800 1536.3500 ;
      RECT 0.0000 1535.9500 1420.0000 1536.0500 ;
      RECT 0.6200 1535.6500 1420.0000 1535.9500 ;
      RECT 0.0000 1532.3500 1420.0000 1535.6500 ;
      RECT 0.0000 1532.0500 1419.3800 1532.3500 ;
      RECT 0.0000 1531.9500 1420.0000 1532.0500 ;
      RECT 0.6200 1531.6500 1420.0000 1531.9500 ;
      RECT 0.0000 1528.3500 1420.0000 1531.6500 ;
      RECT 0.0000 1528.0500 1419.3800 1528.3500 ;
      RECT 0.0000 1527.9500 1420.0000 1528.0500 ;
      RECT 0.6200 1527.6500 1420.0000 1527.9500 ;
      RECT 0.0000 1524.3500 1420.0000 1527.6500 ;
      RECT 0.0000 1524.0500 1419.3800 1524.3500 ;
      RECT 0.0000 1523.9500 1420.0000 1524.0500 ;
      RECT 0.6200 1523.6500 1420.0000 1523.9500 ;
      RECT 0.0000 1520.3500 1420.0000 1523.6500 ;
      RECT 0.0000 1520.0500 1419.3800 1520.3500 ;
      RECT 0.0000 1519.9500 1420.0000 1520.0500 ;
      RECT 0.6200 1519.6500 1420.0000 1519.9500 ;
      RECT 0.0000 1516.3500 1420.0000 1519.6500 ;
      RECT 0.0000 1516.0500 1419.3800 1516.3500 ;
      RECT 0.0000 1515.9500 1420.0000 1516.0500 ;
      RECT 0.6200 1515.6500 1420.0000 1515.9500 ;
      RECT 0.0000 1512.3500 1420.0000 1515.6500 ;
      RECT 0.0000 1512.0500 1419.3800 1512.3500 ;
      RECT 0.0000 1511.9500 1420.0000 1512.0500 ;
      RECT 0.6200 1511.6500 1420.0000 1511.9500 ;
      RECT 0.0000 1508.3500 1420.0000 1511.6500 ;
      RECT 0.0000 1508.0500 1419.3800 1508.3500 ;
      RECT 0.0000 1507.9500 1420.0000 1508.0500 ;
      RECT 0.6200 1507.6500 1420.0000 1507.9500 ;
      RECT 0.0000 1504.3500 1420.0000 1507.6500 ;
      RECT 0.0000 1504.0500 1419.3800 1504.3500 ;
      RECT 0.0000 1503.9500 1420.0000 1504.0500 ;
      RECT 0.6200 1503.6500 1420.0000 1503.9500 ;
      RECT 0.0000 1500.3500 1420.0000 1503.6500 ;
      RECT 0.0000 1500.0500 1419.3800 1500.3500 ;
      RECT 0.0000 1499.9500 1420.0000 1500.0500 ;
      RECT 0.6200 1499.6500 1420.0000 1499.9500 ;
      RECT 0.0000 1496.3500 1420.0000 1499.6500 ;
      RECT 0.0000 1496.0500 1419.3800 1496.3500 ;
      RECT 0.0000 1495.9500 1420.0000 1496.0500 ;
      RECT 0.6200 1495.6500 1420.0000 1495.9500 ;
      RECT 0.0000 1492.3500 1420.0000 1495.6500 ;
      RECT 0.0000 1492.0500 1419.3800 1492.3500 ;
      RECT 0.0000 1491.9500 1420.0000 1492.0500 ;
      RECT 0.6200 1491.6500 1420.0000 1491.9500 ;
      RECT 0.0000 1488.3500 1420.0000 1491.6500 ;
      RECT 0.0000 1488.0500 1419.3800 1488.3500 ;
      RECT 0.0000 1487.9500 1420.0000 1488.0500 ;
      RECT 0.6200 1487.6500 1420.0000 1487.9500 ;
      RECT 0.0000 1484.3500 1420.0000 1487.6500 ;
      RECT 0.0000 1484.0500 1419.3800 1484.3500 ;
      RECT 0.0000 1483.9500 1420.0000 1484.0500 ;
      RECT 0.6200 1483.6500 1420.0000 1483.9500 ;
      RECT 0.0000 1480.3500 1420.0000 1483.6500 ;
      RECT 0.0000 1480.0500 1419.3800 1480.3500 ;
      RECT 0.0000 1479.9500 1420.0000 1480.0500 ;
      RECT 0.6200 1479.6500 1420.0000 1479.9500 ;
      RECT 0.0000 1476.3500 1420.0000 1479.6500 ;
      RECT 0.0000 1476.0500 1419.3800 1476.3500 ;
      RECT 0.0000 1475.9500 1420.0000 1476.0500 ;
      RECT 0.6200 1475.6500 1420.0000 1475.9500 ;
      RECT 0.0000 1472.3500 1420.0000 1475.6500 ;
      RECT 0.0000 1472.0500 1419.3800 1472.3500 ;
      RECT 0.0000 1471.9500 1420.0000 1472.0500 ;
      RECT 0.6200 1471.6500 1420.0000 1471.9500 ;
      RECT 0.0000 1468.3500 1420.0000 1471.6500 ;
      RECT 0.0000 1468.0500 1419.3800 1468.3500 ;
      RECT 0.0000 1467.9500 1420.0000 1468.0500 ;
      RECT 0.6200 1467.6500 1420.0000 1467.9500 ;
      RECT 0.0000 1464.3500 1420.0000 1467.6500 ;
      RECT 0.0000 1464.0500 1419.3800 1464.3500 ;
      RECT 0.0000 1463.9500 1420.0000 1464.0500 ;
      RECT 0.6200 1463.6500 1420.0000 1463.9500 ;
      RECT 0.0000 1460.3500 1420.0000 1463.6500 ;
      RECT 0.0000 1460.0500 1419.3800 1460.3500 ;
      RECT 0.0000 1459.9500 1420.0000 1460.0500 ;
      RECT 0.6200 1459.6500 1420.0000 1459.9500 ;
      RECT 0.0000 1456.3500 1420.0000 1459.6500 ;
      RECT 0.0000 1456.0500 1419.3800 1456.3500 ;
      RECT 0.0000 1455.9500 1420.0000 1456.0500 ;
      RECT 0.6200 1455.6500 1420.0000 1455.9500 ;
      RECT 0.0000 1452.3500 1420.0000 1455.6500 ;
      RECT 0.0000 1452.0500 1419.3800 1452.3500 ;
      RECT 0.0000 1451.9500 1420.0000 1452.0500 ;
      RECT 0.6200 1451.6500 1420.0000 1451.9500 ;
      RECT 0.0000 1449.9500 1420.0000 1451.6500 ;
      RECT 0.6200 1449.6500 1420.0000 1449.9500 ;
      RECT 0.0000 1448.3500 1420.0000 1449.6500 ;
      RECT 0.0000 1448.0500 1419.3800 1448.3500 ;
      RECT 0.0000 1447.9500 1420.0000 1448.0500 ;
      RECT 0.6200 1447.6500 1420.0000 1447.9500 ;
      RECT 0.0000 1445.9500 1420.0000 1447.6500 ;
      RECT 0.6200 1445.6500 1420.0000 1445.9500 ;
      RECT 0.0000 1444.3500 1420.0000 1445.6500 ;
      RECT 0.0000 1444.0500 1419.3800 1444.3500 ;
      RECT 0.0000 1443.9500 1420.0000 1444.0500 ;
      RECT 0.6200 1443.6500 1420.0000 1443.9500 ;
      RECT 0.0000 1441.9500 1420.0000 1443.6500 ;
      RECT 0.6200 1441.6500 1420.0000 1441.9500 ;
      RECT 0.0000 1440.3500 1420.0000 1441.6500 ;
      RECT 0.0000 1440.0500 1419.3800 1440.3500 ;
      RECT 0.0000 1439.9500 1420.0000 1440.0500 ;
      RECT 0.6200 1439.6500 1420.0000 1439.9500 ;
      RECT 0.0000 1437.9500 1420.0000 1439.6500 ;
      RECT 0.6200 1437.6500 1420.0000 1437.9500 ;
      RECT 0.0000 1436.3500 1420.0000 1437.6500 ;
      RECT 0.0000 1436.0500 1419.3800 1436.3500 ;
      RECT 0.0000 1435.9500 1420.0000 1436.0500 ;
      RECT 0.6200 1435.6500 1420.0000 1435.9500 ;
      RECT 0.0000 1433.9500 1420.0000 1435.6500 ;
      RECT 0.6200 1433.6500 1420.0000 1433.9500 ;
      RECT 0.0000 1432.3500 1420.0000 1433.6500 ;
      RECT 0.0000 1432.0500 1419.3800 1432.3500 ;
      RECT 0.0000 1431.9500 1420.0000 1432.0500 ;
      RECT 0.6200 1431.6500 1420.0000 1431.9500 ;
      RECT 0.0000 1429.9500 1420.0000 1431.6500 ;
      RECT 0.6200 1429.6500 1420.0000 1429.9500 ;
      RECT 0.0000 1428.3500 1420.0000 1429.6500 ;
      RECT 0.0000 1428.0500 1419.3800 1428.3500 ;
      RECT 0.0000 1427.9500 1420.0000 1428.0500 ;
      RECT 0.6200 1427.6500 1420.0000 1427.9500 ;
      RECT 0.0000 1425.9500 1420.0000 1427.6500 ;
      RECT 0.6200 1425.6500 1420.0000 1425.9500 ;
      RECT 0.0000 1424.3500 1420.0000 1425.6500 ;
      RECT 0.0000 1424.0500 1419.3800 1424.3500 ;
      RECT 0.0000 1423.9500 1420.0000 1424.0500 ;
      RECT 0.6200 1423.6500 1420.0000 1423.9500 ;
      RECT 0.0000 1421.9500 1420.0000 1423.6500 ;
      RECT 0.6200 1421.6500 1420.0000 1421.9500 ;
      RECT 0.0000 1420.3500 1420.0000 1421.6500 ;
      RECT 0.0000 1420.0500 1419.3800 1420.3500 ;
      RECT 0.0000 1419.9500 1420.0000 1420.0500 ;
      RECT 0.6200 1419.6500 1420.0000 1419.9500 ;
      RECT 0.0000 1417.9500 1420.0000 1419.6500 ;
      RECT 0.6200 1417.6500 1420.0000 1417.9500 ;
      RECT 0.0000 1416.3500 1420.0000 1417.6500 ;
      RECT 0.0000 1416.0500 1419.3800 1416.3500 ;
      RECT 0.0000 1415.9500 1420.0000 1416.0500 ;
      RECT 0.6200 1415.6500 1420.0000 1415.9500 ;
      RECT 0.0000 1413.9500 1420.0000 1415.6500 ;
      RECT 0.6200 1413.6500 1420.0000 1413.9500 ;
      RECT 0.0000 1412.3500 1420.0000 1413.6500 ;
      RECT 0.0000 1412.0500 1419.3800 1412.3500 ;
      RECT 0.0000 1411.9500 1420.0000 1412.0500 ;
      RECT 0.6200 1411.6500 1420.0000 1411.9500 ;
      RECT 0.0000 1409.9500 1420.0000 1411.6500 ;
      RECT 0.6200 1409.6500 1420.0000 1409.9500 ;
      RECT 0.0000 1408.3500 1420.0000 1409.6500 ;
      RECT 0.0000 1408.0500 1419.3800 1408.3500 ;
      RECT 0.0000 1407.9500 1420.0000 1408.0500 ;
      RECT 0.6200 1407.6500 1420.0000 1407.9500 ;
      RECT 0.0000 1405.9500 1420.0000 1407.6500 ;
      RECT 0.6200 1405.6500 1420.0000 1405.9500 ;
      RECT 0.0000 1404.3500 1420.0000 1405.6500 ;
      RECT 0.0000 1404.0500 1419.3800 1404.3500 ;
      RECT 0.0000 1403.9500 1420.0000 1404.0500 ;
      RECT 0.6200 1403.6500 1420.0000 1403.9500 ;
      RECT 0.0000 1401.9500 1420.0000 1403.6500 ;
      RECT 0.6200 1401.6500 1420.0000 1401.9500 ;
      RECT 0.0000 1400.3500 1420.0000 1401.6500 ;
      RECT 0.0000 1400.0500 1419.3800 1400.3500 ;
      RECT 0.0000 1399.9500 1420.0000 1400.0500 ;
      RECT 0.6200 1399.6500 1420.0000 1399.9500 ;
      RECT 0.0000 1397.9500 1420.0000 1399.6500 ;
      RECT 0.6200 1397.6500 1420.0000 1397.9500 ;
      RECT 0.0000 1396.3500 1420.0000 1397.6500 ;
      RECT 0.0000 1396.0500 1419.3800 1396.3500 ;
      RECT 0.0000 1395.9500 1420.0000 1396.0500 ;
      RECT 0.6200 1395.6500 1420.0000 1395.9500 ;
      RECT 0.0000 1393.9500 1420.0000 1395.6500 ;
      RECT 0.6200 1393.6500 1420.0000 1393.9500 ;
      RECT 0.0000 1392.3500 1420.0000 1393.6500 ;
      RECT 0.0000 1392.0500 1419.3800 1392.3500 ;
      RECT 0.0000 1391.9500 1420.0000 1392.0500 ;
      RECT 0.6200 1391.6500 1420.0000 1391.9500 ;
      RECT 0.0000 1389.9500 1420.0000 1391.6500 ;
      RECT 0.6200 1389.6500 1420.0000 1389.9500 ;
      RECT 0.0000 1388.3500 1420.0000 1389.6500 ;
      RECT 0.0000 1388.0500 1419.3800 1388.3500 ;
      RECT 0.0000 1387.9500 1420.0000 1388.0500 ;
      RECT 0.6200 1387.6500 1420.0000 1387.9500 ;
      RECT 0.0000 1385.9500 1420.0000 1387.6500 ;
      RECT 0.6200 1385.6500 1420.0000 1385.9500 ;
      RECT 0.0000 1384.3500 1420.0000 1385.6500 ;
      RECT 0.0000 1384.0500 1419.3800 1384.3500 ;
      RECT 0.0000 1383.9500 1420.0000 1384.0500 ;
      RECT 0.6200 1383.6500 1420.0000 1383.9500 ;
      RECT 0.0000 1381.9500 1420.0000 1383.6500 ;
      RECT 0.6200 1381.6500 1420.0000 1381.9500 ;
      RECT 0.0000 1380.3500 1420.0000 1381.6500 ;
      RECT 0.0000 1380.0500 1419.3800 1380.3500 ;
      RECT 0.0000 1379.9500 1420.0000 1380.0500 ;
      RECT 0.6200 1379.6500 1420.0000 1379.9500 ;
      RECT 0.0000 1377.9500 1420.0000 1379.6500 ;
      RECT 0.6200 1377.6500 1420.0000 1377.9500 ;
      RECT 0.0000 1376.3500 1420.0000 1377.6500 ;
      RECT 0.0000 1376.0500 1419.3800 1376.3500 ;
      RECT 0.0000 1375.9500 1420.0000 1376.0500 ;
      RECT 0.6200 1375.6500 1420.0000 1375.9500 ;
      RECT 0.0000 1373.9500 1420.0000 1375.6500 ;
      RECT 0.6200 1373.6500 1420.0000 1373.9500 ;
      RECT 0.0000 1372.3500 1420.0000 1373.6500 ;
      RECT 0.0000 1372.0500 1419.3800 1372.3500 ;
      RECT 0.0000 1371.9500 1420.0000 1372.0500 ;
      RECT 0.6200 1371.6500 1420.0000 1371.9500 ;
      RECT 0.0000 1369.9500 1420.0000 1371.6500 ;
      RECT 0.6200 1369.6500 1420.0000 1369.9500 ;
      RECT 0.0000 1368.3500 1420.0000 1369.6500 ;
      RECT 0.0000 1368.0500 1419.3800 1368.3500 ;
      RECT 0.0000 1367.9500 1420.0000 1368.0500 ;
      RECT 0.6200 1367.6500 1420.0000 1367.9500 ;
      RECT 0.0000 1364.3500 1420.0000 1367.6500 ;
      RECT 0.0000 1364.0500 1419.3800 1364.3500 ;
      RECT 0.0000 1363.9500 1420.0000 1364.0500 ;
      RECT 0.6200 1363.6500 1420.0000 1363.9500 ;
      RECT 0.0000 1360.3500 1420.0000 1363.6500 ;
      RECT 0.0000 1360.0500 1419.3800 1360.3500 ;
      RECT 0.0000 1359.9500 1420.0000 1360.0500 ;
      RECT 0.6200 1359.6500 1420.0000 1359.9500 ;
      RECT 0.0000 1356.3500 1420.0000 1359.6500 ;
      RECT 0.0000 1356.0500 1419.3800 1356.3500 ;
      RECT 0.0000 1355.9500 1420.0000 1356.0500 ;
      RECT 0.6200 1355.6500 1420.0000 1355.9500 ;
      RECT 0.0000 1352.3500 1420.0000 1355.6500 ;
      RECT 0.0000 1352.0500 1419.3800 1352.3500 ;
      RECT 0.0000 1351.9500 1420.0000 1352.0500 ;
      RECT 0.6200 1351.6500 1420.0000 1351.9500 ;
      RECT 0.0000 1348.3500 1420.0000 1351.6500 ;
      RECT 0.0000 1348.0500 1419.3800 1348.3500 ;
      RECT 0.0000 1347.9500 1420.0000 1348.0500 ;
      RECT 0.6200 1347.6500 1420.0000 1347.9500 ;
      RECT 0.0000 1344.3500 1420.0000 1347.6500 ;
      RECT 0.0000 1344.0500 1419.3800 1344.3500 ;
      RECT 0.0000 1343.9500 1420.0000 1344.0500 ;
      RECT 0.6200 1343.6500 1420.0000 1343.9500 ;
      RECT 0.0000 1340.3500 1420.0000 1343.6500 ;
      RECT 0.0000 1340.0500 1419.3800 1340.3500 ;
      RECT 0.0000 1339.9500 1420.0000 1340.0500 ;
      RECT 0.6200 1339.6500 1420.0000 1339.9500 ;
      RECT 0.0000 1336.3500 1420.0000 1339.6500 ;
      RECT 0.0000 1336.0500 1419.3800 1336.3500 ;
      RECT 0.0000 1335.9500 1420.0000 1336.0500 ;
      RECT 0.6200 1335.6500 1420.0000 1335.9500 ;
      RECT 0.0000 1332.3500 1420.0000 1335.6500 ;
      RECT 0.0000 1332.0500 1419.3800 1332.3500 ;
      RECT 0.0000 1331.9500 1420.0000 1332.0500 ;
      RECT 0.6200 1331.6500 1420.0000 1331.9500 ;
      RECT 0.0000 1328.3500 1420.0000 1331.6500 ;
      RECT 0.0000 1328.0500 1419.3800 1328.3500 ;
      RECT 0.0000 1327.9500 1420.0000 1328.0500 ;
      RECT 0.6200 1327.6500 1420.0000 1327.9500 ;
      RECT 0.0000 1324.3500 1420.0000 1327.6500 ;
      RECT 0.0000 1324.0500 1419.3800 1324.3500 ;
      RECT 0.0000 1323.9500 1420.0000 1324.0500 ;
      RECT 0.6200 1323.6500 1420.0000 1323.9500 ;
      RECT 0.0000 1320.3500 1420.0000 1323.6500 ;
      RECT 0.0000 1320.0500 1419.3800 1320.3500 ;
      RECT 0.0000 1319.9500 1420.0000 1320.0500 ;
      RECT 0.6200 1319.6500 1420.0000 1319.9500 ;
      RECT 0.0000 1316.3500 1420.0000 1319.6500 ;
      RECT 0.0000 1316.0500 1419.3800 1316.3500 ;
      RECT 0.0000 1315.9500 1420.0000 1316.0500 ;
      RECT 0.6200 1315.6500 1420.0000 1315.9500 ;
      RECT 0.0000 1312.3500 1420.0000 1315.6500 ;
      RECT 0.0000 1312.0500 1419.3800 1312.3500 ;
      RECT 0.0000 1311.9500 1420.0000 1312.0500 ;
      RECT 0.6200 1311.6500 1420.0000 1311.9500 ;
      RECT 0.0000 1308.3500 1420.0000 1311.6500 ;
      RECT 0.0000 1308.0500 1419.3800 1308.3500 ;
      RECT 0.0000 1307.9500 1420.0000 1308.0500 ;
      RECT 0.6200 1307.6500 1420.0000 1307.9500 ;
      RECT 0.0000 1304.3500 1420.0000 1307.6500 ;
      RECT 0.0000 1304.0500 1419.3800 1304.3500 ;
      RECT 0.0000 1303.9500 1420.0000 1304.0500 ;
      RECT 0.6200 1303.6500 1420.0000 1303.9500 ;
      RECT 0.0000 1300.3500 1420.0000 1303.6500 ;
      RECT 0.0000 1300.0500 1419.3800 1300.3500 ;
      RECT 0.0000 1299.9500 1420.0000 1300.0500 ;
      RECT 0.6200 1299.6500 1420.0000 1299.9500 ;
      RECT 0.0000 1296.3500 1420.0000 1299.6500 ;
      RECT 0.0000 1296.0500 1419.3800 1296.3500 ;
      RECT 0.0000 1295.9500 1420.0000 1296.0500 ;
      RECT 0.6200 1295.6500 1420.0000 1295.9500 ;
      RECT 0.0000 1292.3500 1420.0000 1295.6500 ;
      RECT 0.0000 1292.0500 1419.3800 1292.3500 ;
      RECT 0.0000 1291.9500 1420.0000 1292.0500 ;
      RECT 0.6200 1291.6500 1420.0000 1291.9500 ;
      RECT 0.0000 1288.3500 1420.0000 1291.6500 ;
      RECT 0.0000 1288.0500 1419.3800 1288.3500 ;
      RECT 0.0000 1287.9500 1420.0000 1288.0500 ;
      RECT 0.6200 1287.6500 1420.0000 1287.9500 ;
      RECT 0.0000 1284.3500 1420.0000 1287.6500 ;
      RECT 0.0000 1284.0500 1419.3800 1284.3500 ;
      RECT 0.0000 1283.9500 1420.0000 1284.0500 ;
      RECT 0.6200 1283.6500 1420.0000 1283.9500 ;
      RECT 0.0000 1280.3500 1420.0000 1283.6500 ;
      RECT 0.0000 1280.0500 1419.3800 1280.3500 ;
      RECT 0.0000 1279.9500 1420.0000 1280.0500 ;
      RECT 0.6200 1279.6500 1420.0000 1279.9500 ;
      RECT 0.0000 1276.3500 1420.0000 1279.6500 ;
      RECT 0.0000 1276.0500 1419.3800 1276.3500 ;
      RECT 0.0000 1275.9500 1420.0000 1276.0500 ;
      RECT 0.6200 1275.6500 1420.0000 1275.9500 ;
      RECT 0.0000 1272.3500 1420.0000 1275.6500 ;
      RECT 0.0000 1272.0500 1419.3800 1272.3500 ;
      RECT 0.0000 1271.9500 1420.0000 1272.0500 ;
      RECT 0.6200 1271.6500 1420.0000 1271.9500 ;
      RECT 0.0000 1268.3500 1420.0000 1271.6500 ;
      RECT 0.0000 1268.0500 1419.3800 1268.3500 ;
      RECT 0.0000 1267.9500 1420.0000 1268.0500 ;
      RECT 0.6200 1267.6500 1420.0000 1267.9500 ;
      RECT 0.0000 1264.3500 1420.0000 1267.6500 ;
      RECT 0.0000 1264.0500 1419.3800 1264.3500 ;
      RECT 0.0000 1263.9500 1420.0000 1264.0500 ;
      RECT 0.6200 1263.6500 1420.0000 1263.9500 ;
      RECT 0.0000 1260.3500 1420.0000 1263.6500 ;
      RECT 0.0000 1260.0500 1419.3800 1260.3500 ;
      RECT 0.0000 1259.9500 1420.0000 1260.0500 ;
      RECT 0.6200 1259.6500 1420.0000 1259.9500 ;
      RECT 0.0000 1256.3500 1420.0000 1259.6500 ;
      RECT 0.0000 1256.0500 1419.3800 1256.3500 ;
      RECT 0.0000 1255.9500 1420.0000 1256.0500 ;
      RECT 0.6200 1255.6500 1420.0000 1255.9500 ;
      RECT 0.0000 1252.3500 1420.0000 1255.6500 ;
      RECT 0.0000 1252.0500 1419.3800 1252.3500 ;
      RECT 0.0000 1251.9500 1420.0000 1252.0500 ;
      RECT 0.6200 1251.6500 1420.0000 1251.9500 ;
      RECT 0.0000 1248.3500 1420.0000 1251.6500 ;
      RECT 0.0000 1248.0500 1419.3800 1248.3500 ;
      RECT 0.0000 1247.9500 1420.0000 1248.0500 ;
      RECT 0.6200 1247.6500 1420.0000 1247.9500 ;
      RECT 0.0000 1244.3500 1420.0000 1247.6500 ;
      RECT 0.0000 1244.0500 1419.3800 1244.3500 ;
      RECT 0.0000 1243.9500 1420.0000 1244.0500 ;
      RECT 0.6200 1243.6500 1420.0000 1243.9500 ;
      RECT 0.0000 1240.3500 1420.0000 1243.6500 ;
      RECT 0.0000 1240.0500 1419.3800 1240.3500 ;
      RECT 0.0000 1239.9500 1420.0000 1240.0500 ;
      RECT 0.6200 1239.6500 1420.0000 1239.9500 ;
      RECT 0.0000 1236.3500 1420.0000 1239.6500 ;
      RECT 0.0000 1236.0500 1419.3800 1236.3500 ;
      RECT 0.0000 1235.9500 1420.0000 1236.0500 ;
      RECT 0.6200 1235.6500 1420.0000 1235.9500 ;
      RECT 0.0000 1232.3500 1420.0000 1235.6500 ;
      RECT 0.0000 1232.0500 1419.3800 1232.3500 ;
      RECT 0.0000 1231.9500 1420.0000 1232.0500 ;
      RECT 0.6200 1231.6500 1420.0000 1231.9500 ;
      RECT 0.0000 1228.3500 1420.0000 1231.6500 ;
      RECT 0.0000 1228.0500 1419.3800 1228.3500 ;
      RECT 0.0000 1227.9500 1420.0000 1228.0500 ;
      RECT 0.6200 1227.6500 1420.0000 1227.9500 ;
      RECT 0.0000 1224.3500 1420.0000 1227.6500 ;
      RECT 0.0000 1224.0500 1419.3800 1224.3500 ;
      RECT 0.0000 1223.9500 1420.0000 1224.0500 ;
      RECT 0.6200 1223.6500 1420.0000 1223.9500 ;
      RECT 0.0000 1220.3500 1420.0000 1223.6500 ;
      RECT 0.0000 1220.0500 1419.3800 1220.3500 ;
      RECT 0.0000 1219.9500 1420.0000 1220.0500 ;
      RECT 0.6200 1219.6500 1420.0000 1219.9500 ;
      RECT 0.0000 1216.3500 1420.0000 1219.6500 ;
      RECT 0.0000 1216.0500 1419.3800 1216.3500 ;
      RECT 0.0000 1215.9500 1420.0000 1216.0500 ;
      RECT 0.6200 1215.6500 1420.0000 1215.9500 ;
      RECT 0.0000 1212.3500 1420.0000 1215.6500 ;
      RECT 0.0000 1212.0500 1419.3800 1212.3500 ;
      RECT 0.0000 1211.9500 1420.0000 1212.0500 ;
      RECT 0.6200 1211.6500 1420.0000 1211.9500 ;
      RECT 0.0000 1208.3500 1420.0000 1211.6500 ;
      RECT 0.0000 1208.0500 1419.3800 1208.3500 ;
      RECT 0.0000 1207.9500 1420.0000 1208.0500 ;
      RECT 0.6200 1207.6500 1420.0000 1207.9500 ;
      RECT 0.0000 1204.3500 1420.0000 1207.6500 ;
      RECT 0.0000 1204.0500 1419.3800 1204.3500 ;
      RECT 0.0000 1203.9500 1420.0000 1204.0500 ;
      RECT 0.6200 1203.6500 1420.0000 1203.9500 ;
      RECT 0.0000 1200.3500 1420.0000 1203.6500 ;
      RECT 0.0000 1200.0500 1419.3800 1200.3500 ;
      RECT 0.0000 1199.9500 1420.0000 1200.0500 ;
      RECT 0.6200 1199.6500 1420.0000 1199.9500 ;
      RECT 0.0000 1196.3500 1420.0000 1199.6500 ;
      RECT 0.0000 1196.0500 1419.3800 1196.3500 ;
      RECT 0.0000 1195.9500 1420.0000 1196.0500 ;
      RECT 0.6200 1195.6500 1420.0000 1195.9500 ;
      RECT 0.0000 1192.3500 1420.0000 1195.6500 ;
      RECT 0.0000 1192.0500 1419.3800 1192.3500 ;
      RECT 0.0000 1191.9500 1420.0000 1192.0500 ;
      RECT 0.6200 1191.6500 1420.0000 1191.9500 ;
      RECT 0.0000 1188.3500 1420.0000 1191.6500 ;
      RECT 0.0000 1188.0500 1419.3800 1188.3500 ;
      RECT 0.0000 1187.9500 1420.0000 1188.0500 ;
      RECT 0.6200 1187.6500 1420.0000 1187.9500 ;
      RECT 0.0000 1184.3500 1420.0000 1187.6500 ;
      RECT 0.0000 1184.0500 1419.3800 1184.3500 ;
      RECT 0.0000 1183.9500 1420.0000 1184.0500 ;
      RECT 0.6200 1183.6500 1420.0000 1183.9500 ;
      RECT 0.0000 1180.3500 1420.0000 1183.6500 ;
      RECT 0.0000 1180.0500 1419.3800 1180.3500 ;
      RECT 0.0000 1179.9500 1420.0000 1180.0500 ;
      RECT 0.6200 1179.6500 1420.0000 1179.9500 ;
      RECT 0.0000 1176.3500 1420.0000 1179.6500 ;
      RECT 0.0000 1176.0500 1419.3800 1176.3500 ;
      RECT 0.0000 1175.9500 1420.0000 1176.0500 ;
      RECT 0.6200 1175.6500 1420.0000 1175.9500 ;
      RECT 0.0000 1172.3500 1420.0000 1175.6500 ;
      RECT 0.0000 1172.0500 1419.3800 1172.3500 ;
      RECT 0.0000 1171.9500 1420.0000 1172.0500 ;
      RECT 0.6200 1171.6500 1420.0000 1171.9500 ;
      RECT 0.0000 1168.3500 1420.0000 1171.6500 ;
      RECT 0.0000 1168.0500 1419.3800 1168.3500 ;
      RECT 0.0000 1167.9500 1420.0000 1168.0500 ;
      RECT 0.6200 1167.6500 1420.0000 1167.9500 ;
      RECT 0.0000 1164.3500 1420.0000 1167.6500 ;
      RECT 0.0000 1164.0500 1419.3800 1164.3500 ;
      RECT 0.0000 1163.9500 1420.0000 1164.0500 ;
      RECT 0.6200 1163.6500 1420.0000 1163.9500 ;
      RECT 0.0000 1160.3500 1420.0000 1163.6500 ;
      RECT 0.0000 1160.0500 1419.3800 1160.3500 ;
      RECT 0.0000 1159.9500 1420.0000 1160.0500 ;
      RECT 0.6200 1159.6500 1420.0000 1159.9500 ;
      RECT 0.0000 1156.3500 1420.0000 1159.6500 ;
      RECT 0.0000 1156.0500 1419.3800 1156.3500 ;
      RECT 0.0000 1155.9500 1420.0000 1156.0500 ;
      RECT 0.6200 1155.6500 1420.0000 1155.9500 ;
      RECT 0.0000 1152.3500 1420.0000 1155.6500 ;
      RECT 0.0000 1152.0500 1419.3800 1152.3500 ;
      RECT 0.0000 1148.3500 1420.0000 1152.0500 ;
      RECT 0.0000 1148.0500 1419.3800 1148.3500 ;
      RECT 0.0000 1144.3500 1420.0000 1148.0500 ;
      RECT 0.0000 1144.0500 1419.3800 1144.3500 ;
      RECT 0.0000 1140.3500 1420.0000 1144.0500 ;
      RECT 0.0000 1140.0500 1419.3800 1140.3500 ;
      RECT 0.0000 1136.3500 1420.0000 1140.0500 ;
      RECT 0.0000 1136.0500 1419.3800 1136.3500 ;
      RECT 0.0000 1132.3500 1420.0000 1136.0500 ;
      RECT 0.0000 1132.0500 1419.3800 1132.3500 ;
      RECT 0.0000 1128.3500 1420.0000 1132.0500 ;
      RECT 0.0000 1128.0500 1419.3800 1128.3500 ;
      RECT 0.0000 1124.3500 1420.0000 1128.0500 ;
      RECT 0.0000 1124.0500 1419.3800 1124.3500 ;
      RECT 0.0000 1120.3500 1420.0000 1124.0500 ;
      RECT 0.0000 1120.0500 1419.3800 1120.3500 ;
      RECT 0.0000 1116.3500 1420.0000 1120.0500 ;
      RECT 0.0000 1116.0500 1419.3800 1116.3500 ;
      RECT 0.0000 1112.3500 1420.0000 1116.0500 ;
      RECT 0.0000 1112.0500 1419.3800 1112.3500 ;
      RECT 0.0000 1108.3500 1420.0000 1112.0500 ;
      RECT 0.0000 1108.0500 1419.3800 1108.3500 ;
      RECT 0.0000 1104.3500 1420.0000 1108.0500 ;
      RECT 0.0000 1104.0500 1419.3800 1104.3500 ;
      RECT 0.0000 1100.3500 1420.0000 1104.0500 ;
      RECT 0.0000 1100.0500 1419.3800 1100.3500 ;
      RECT 0.0000 1096.3500 1420.0000 1100.0500 ;
      RECT 0.0000 1096.0500 1419.3800 1096.3500 ;
      RECT 0.0000 1092.3500 1420.0000 1096.0500 ;
      RECT 0.0000 1092.0500 1419.3800 1092.3500 ;
      RECT 0.0000 1088.3500 1420.0000 1092.0500 ;
      RECT 0.0000 1088.0500 1419.3800 1088.3500 ;
      RECT 0.0000 1084.3500 1420.0000 1088.0500 ;
      RECT 0.0000 1084.0500 1419.3800 1084.3500 ;
      RECT 0.0000 1080.3500 1420.0000 1084.0500 ;
      RECT 0.0000 1080.0500 1419.3800 1080.3500 ;
      RECT 0.0000 1076.3500 1420.0000 1080.0500 ;
      RECT 0.0000 1076.0500 1419.3800 1076.3500 ;
      RECT 0.0000 1072.3500 1420.0000 1076.0500 ;
      RECT 0.0000 1072.0500 1419.3800 1072.3500 ;
      RECT 0.0000 1068.3500 1420.0000 1072.0500 ;
      RECT 0.0000 1068.0500 1419.3800 1068.3500 ;
      RECT 0.0000 1064.3500 1420.0000 1068.0500 ;
      RECT 0.0000 1064.0500 1419.3800 1064.3500 ;
      RECT 0.0000 1060.3500 1420.0000 1064.0500 ;
      RECT 0.0000 1060.0500 1419.3800 1060.3500 ;
      RECT 0.0000 1056.3500 1420.0000 1060.0500 ;
      RECT 0.0000 1056.0500 1419.3800 1056.3500 ;
      RECT 0.0000 1052.3500 1420.0000 1056.0500 ;
      RECT 0.0000 1052.0500 1419.3800 1052.3500 ;
      RECT 0.0000 1048.3500 1420.0000 1052.0500 ;
      RECT 0.0000 1048.0500 1419.3800 1048.3500 ;
      RECT 0.0000 1044.3500 1420.0000 1048.0500 ;
      RECT 0.0000 1044.0500 1419.3800 1044.3500 ;
      RECT 0.0000 1040.3500 1420.0000 1044.0500 ;
      RECT 0.0000 1040.0500 1419.3800 1040.3500 ;
      RECT 0.0000 1036.3500 1420.0000 1040.0500 ;
      RECT 0.0000 1036.0500 1419.3800 1036.3500 ;
      RECT 0.0000 1032.3500 1420.0000 1036.0500 ;
      RECT 0.0000 1032.0500 1419.3800 1032.3500 ;
      RECT 0.0000 1028.3500 1420.0000 1032.0500 ;
      RECT 0.0000 1028.0500 1419.3800 1028.3500 ;
      RECT 0.0000 1024.3500 1420.0000 1028.0500 ;
      RECT 0.0000 1024.0500 1419.3800 1024.3500 ;
      RECT 0.0000 1020.3500 1420.0000 1024.0500 ;
      RECT 0.0000 1020.0500 1419.3800 1020.3500 ;
      RECT 0.0000 1016.3500 1420.0000 1020.0500 ;
      RECT 0.0000 1016.0500 1419.3800 1016.3500 ;
      RECT 0.0000 1012.3500 1420.0000 1016.0500 ;
      RECT 0.0000 1012.0500 1419.3800 1012.3500 ;
      RECT 0.0000 1008.3500 1420.0000 1012.0500 ;
      RECT 0.0000 1008.0500 1419.3800 1008.3500 ;
      RECT 0.0000 1004.3500 1420.0000 1008.0500 ;
      RECT 0.0000 1004.0500 1419.3800 1004.3500 ;
      RECT 0.0000 1000.3500 1420.0000 1004.0500 ;
      RECT 0.0000 1000.0500 1419.3800 1000.3500 ;
      RECT 0.0000 996.3500 1420.0000 1000.0500 ;
      RECT 0.0000 996.0500 1419.3800 996.3500 ;
      RECT 0.0000 992.3500 1420.0000 996.0500 ;
      RECT 0.0000 992.0500 1419.3800 992.3500 ;
      RECT 0.0000 988.3500 1420.0000 992.0500 ;
      RECT 0.0000 988.0500 1419.3800 988.3500 ;
      RECT 0.0000 984.3500 1420.0000 988.0500 ;
      RECT 0.0000 984.0500 1419.3800 984.3500 ;
      RECT 0.0000 980.3500 1420.0000 984.0500 ;
      RECT 0.0000 980.0500 1419.3800 980.3500 ;
      RECT 0.0000 976.3500 1420.0000 980.0500 ;
      RECT 0.0000 976.0500 1419.3800 976.3500 ;
      RECT 0.0000 972.3500 1420.0000 976.0500 ;
      RECT 0.0000 972.0500 1419.3800 972.3500 ;
      RECT 0.0000 968.3500 1420.0000 972.0500 ;
      RECT 0.0000 968.0500 1419.3800 968.3500 ;
      RECT 0.0000 964.3500 1420.0000 968.0500 ;
      RECT 0.0000 964.0500 1419.3800 964.3500 ;
      RECT 0.0000 960.3500 1420.0000 964.0500 ;
      RECT 0.0000 960.0500 1419.3800 960.3500 ;
      RECT 0.0000 956.3500 1420.0000 960.0500 ;
      RECT 0.0000 956.0500 1419.3800 956.3500 ;
      RECT 0.0000 952.3500 1420.0000 956.0500 ;
      RECT 0.0000 952.0500 1419.3800 952.3500 ;
      RECT 0.0000 948.3500 1420.0000 952.0500 ;
      RECT 0.0000 948.0500 1419.3800 948.3500 ;
      RECT 0.0000 944.3500 1420.0000 948.0500 ;
      RECT 0.0000 944.0500 1419.3800 944.3500 ;
      RECT 0.0000 940.3500 1420.0000 944.0500 ;
      RECT 0.0000 940.0500 1419.3800 940.3500 ;
      RECT 0.0000 936.3500 1420.0000 940.0500 ;
      RECT 0.0000 936.0500 1419.3800 936.3500 ;
      RECT 0.0000 932.3500 1420.0000 936.0500 ;
      RECT 0.0000 932.0500 1419.3800 932.3500 ;
      RECT 0.0000 928.3500 1420.0000 932.0500 ;
      RECT 0.0000 928.0500 1419.3800 928.3500 ;
      RECT 0.0000 924.3500 1420.0000 928.0500 ;
      RECT 0.0000 924.0500 1419.3800 924.3500 ;
      RECT 0.0000 920.3500 1420.0000 924.0500 ;
      RECT 0.0000 920.0500 1419.3800 920.3500 ;
      RECT 0.0000 916.3500 1420.0000 920.0500 ;
      RECT 0.0000 916.0500 1419.3800 916.3500 ;
      RECT 0.0000 912.3500 1420.0000 916.0500 ;
      RECT 0.0000 912.0500 1419.3800 912.3500 ;
      RECT 0.0000 908.3500 1420.0000 912.0500 ;
      RECT 0.0000 908.0500 1419.3800 908.3500 ;
      RECT 0.0000 904.3500 1420.0000 908.0500 ;
      RECT 0.0000 904.0500 1419.3800 904.3500 ;
      RECT 0.0000 900.3500 1420.0000 904.0500 ;
      RECT 0.0000 900.0500 1419.3800 900.3500 ;
      RECT 0.0000 896.3500 1420.0000 900.0500 ;
      RECT 0.0000 896.0500 1419.3800 896.3500 ;
      RECT 0.0000 892.3500 1420.0000 896.0500 ;
      RECT 0.0000 892.0500 1419.3800 892.3500 ;
      RECT 0.0000 888.3500 1420.0000 892.0500 ;
      RECT 0.0000 888.0500 1419.3800 888.3500 ;
      RECT 0.0000 884.3500 1420.0000 888.0500 ;
      RECT 0.0000 884.0500 1419.3800 884.3500 ;
      RECT 0.0000 880.3500 1420.0000 884.0500 ;
      RECT 0.0000 880.0500 1419.3800 880.3500 ;
      RECT 0.0000 876.3500 1420.0000 880.0500 ;
      RECT 0.0000 876.0500 1419.3800 876.3500 ;
      RECT 0.0000 872.3500 1420.0000 876.0500 ;
      RECT 0.0000 872.0500 1419.3800 872.3500 ;
      RECT 0.0000 868.3500 1420.0000 872.0500 ;
      RECT 0.0000 868.0500 1419.3800 868.3500 ;
      RECT 0.0000 864.3500 1420.0000 868.0500 ;
      RECT 0.0000 864.0500 1419.3800 864.3500 ;
      RECT 0.0000 860.3500 1420.0000 864.0500 ;
      RECT 0.0000 860.0500 1419.3800 860.3500 ;
      RECT 0.0000 856.3500 1420.0000 860.0500 ;
      RECT 0.0000 856.0500 1419.3800 856.3500 ;
      RECT 0.0000 852.3500 1420.0000 856.0500 ;
      RECT 0.0000 852.0500 1419.3800 852.3500 ;
      RECT 0.0000 848.3500 1420.0000 852.0500 ;
      RECT 0.0000 848.0500 1419.3800 848.3500 ;
      RECT 0.0000 844.3500 1420.0000 848.0500 ;
      RECT 0.0000 844.0500 1419.3800 844.3500 ;
      RECT 0.0000 840.3500 1420.0000 844.0500 ;
      RECT 0.0000 840.0500 1419.3800 840.3500 ;
      RECT 0.0000 836.3500 1420.0000 840.0500 ;
      RECT 0.0000 836.0500 1419.3800 836.3500 ;
      RECT 0.0000 832.3500 1420.0000 836.0500 ;
      RECT 0.0000 832.0500 1419.3800 832.3500 ;
      RECT 0.0000 828.3500 1420.0000 832.0500 ;
      RECT 0.0000 828.0500 1419.3800 828.3500 ;
      RECT 0.0000 824.3500 1420.0000 828.0500 ;
      RECT 0.0000 824.0500 1419.3800 824.3500 ;
      RECT 0.0000 820.3500 1420.0000 824.0500 ;
      RECT 0.0000 820.0500 1419.3800 820.3500 ;
      RECT 0.0000 816.3500 1420.0000 820.0500 ;
      RECT 0.0000 816.0500 1419.3800 816.3500 ;
      RECT 0.0000 812.3500 1420.0000 816.0500 ;
      RECT 0.0000 812.0500 1419.3800 812.3500 ;
      RECT 0.0000 808.3500 1420.0000 812.0500 ;
      RECT 0.0000 808.0500 1419.3800 808.3500 ;
      RECT 0.0000 804.3500 1420.0000 808.0500 ;
      RECT 0.0000 804.0500 1419.3800 804.3500 ;
      RECT 0.0000 800.3500 1420.0000 804.0500 ;
      RECT 0.0000 800.0500 1419.3800 800.3500 ;
      RECT 0.0000 796.3500 1420.0000 800.0500 ;
      RECT 0.0000 796.0500 1419.3800 796.3500 ;
      RECT 0.0000 792.3500 1420.0000 796.0500 ;
      RECT 0.0000 792.0500 1419.3800 792.3500 ;
      RECT 0.0000 788.3500 1420.0000 792.0500 ;
      RECT 0.0000 788.0500 1419.3800 788.3500 ;
      RECT 0.0000 784.3500 1420.0000 788.0500 ;
      RECT 0.0000 784.0500 1419.3800 784.3500 ;
      RECT 0.0000 780.3500 1420.0000 784.0500 ;
      RECT 0.0000 780.0500 1419.3800 780.3500 ;
      RECT 0.0000 776.3500 1420.0000 780.0500 ;
      RECT 0.0000 776.0500 1419.3800 776.3500 ;
      RECT 0.0000 772.3500 1420.0000 776.0500 ;
      RECT 0.0000 772.0500 1419.3800 772.3500 ;
      RECT 0.0000 0.0000 1420.0000 772.0500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
  END
END fullchip

END LIBRARY
