##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 18:15:56 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 1120.0000 BY 1120.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 591.7500 0.5200 591.8500 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 685.8500 0.0000 685.9500 0.5200 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 681.8500 0.0000 681.9500 0.5200 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 677.8500 0.0000 677.9500 0.5200 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 673.8500 0.0000 673.9500 0.5200 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 669.8500 0.0000 669.9500 0.5200 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.8500 0.0000 665.9500 0.5200 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 661.8500 0.0000 661.9500 0.5200 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 657.8500 0.0000 657.9500 0.5200 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 653.8500 0.0000 653.9500 0.5200 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 649.8500 0.0000 649.9500 0.5200 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 645.8500 0.0000 645.9500 0.5200 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 641.8500 0.0000 641.9500 0.5200 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 637.8500 0.0000 637.9500 0.5200 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 633.8500 0.0000 633.9500 0.5200 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 629.8500 0.0000 629.9500 0.5200 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 625.8500 0.0000 625.9500 0.5200 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 621.8500 0.0000 621.9500 0.5200 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 617.8500 0.0000 617.9500 0.5200 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 613.8500 0.0000 613.9500 0.5200 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 609.8500 0.0000 609.9500 0.5200 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 605.8500 0.0000 605.9500 0.5200 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 601.8500 0.0000 601.9500 0.5200 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 597.8500 0.0000 597.9500 0.5200 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 593.8500 0.0000 593.9500 0.5200 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 589.8500 0.0000 589.9500 0.5200 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 585.8500 0.0000 585.9500 0.5200 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 581.8500 0.0000 581.9500 0.5200 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 577.8500 0.0000 577.9500 0.5200 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 573.8500 0.0000 573.9500 0.5200 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 569.8500 0.0000 569.9500 0.5200 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 565.8500 0.0000 565.9500 0.5200 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 561.8500 0.0000 561.9500 0.5200 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 557.8500 0.0000 557.9500 0.5200 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 553.8500 0.0000 553.9500 0.5200 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 549.8500 0.0000 549.9500 0.5200 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 545.8500 0.0000 545.9500 0.5200 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 541.8500 0.0000 541.9500 0.5200 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 537.8500 0.0000 537.9500 0.5200 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 533.8500 0.0000 533.9500 0.5200 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 529.8500 0.0000 529.9500 0.5200 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 525.8500 0.0000 525.9500 0.5200 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 521.8500 0.0000 521.9500 0.5200 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 517.8500 0.0000 517.9500 0.5200 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 513.8500 0.0000 513.9500 0.5200 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 509.8500 0.0000 509.9500 0.5200 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 505.8500 0.0000 505.9500 0.5200 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 501.8500 0.0000 501.9500 0.5200 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 497.8500 0.0000 497.9500 0.5200 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 493.8500 0.0000 493.9500 0.5200 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 489.8500 0.0000 489.9500 0.5200 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 485.8500 0.0000 485.9500 0.5200 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 481.8500 0.0000 481.9500 0.5200 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 477.8500 0.0000 477.9500 0.5200 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 473.8500 0.0000 473.9500 0.5200 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 469.8500 0.0000 469.9500 0.5200 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 465.8500 0.0000 465.9500 0.5200 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 461.8500 0.0000 461.9500 0.5200 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.8500 0.0000 457.9500 0.5200 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 453.8500 0.0000 453.9500 0.5200 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.8500 0.0000 449.9500 0.5200 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.8500 0.0000 445.9500 0.5200 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.8500 0.0000 441.9500 0.5200 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 437.8500 0.0000 437.9500 0.5200 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.8500 0.0000 433.9500 0.5200 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 877.8500 1119.4800 877.9500 1120.0000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 873.8500 1119.4800 873.9500 1120.0000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 869.8500 1119.4800 869.9500 1120.0000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 865.8500 1119.4800 865.9500 1120.0000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 861.8500 1119.4800 861.9500 1120.0000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 857.8500 1119.4800 857.9500 1120.0000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 853.8500 1119.4800 853.9500 1120.0000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 849.8500 1119.4800 849.9500 1120.0000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 845.8500 1119.4800 845.9500 1120.0000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 841.8500 1119.4800 841.9500 1120.0000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 837.8500 1119.4800 837.9500 1120.0000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 833.8500 1119.4800 833.9500 1120.0000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 829.8500 1119.4800 829.9500 1120.0000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 825.8500 1119.4800 825.9500 1120.0000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 821.8500 1119.4800 821.9500 1120.0000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 817.8500 1119.4800 817.9500 1120.0000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 813.8500 1119.4800 813.9500 1120.0000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 809.8500 1119.4800 809.9500 1120.0000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 805.8500 1119.4800 805.9500 1120.0000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 801.8500 1119.4800 801.9500 1120.0000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 797.8500 1119.4800 797.9500 1120.0000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 793.8500 1119.4800 793.9500 1120.0000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 789.8500 1119.4800 789.9500 1120.0000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 785.8500 1119.4800 785.9500 1120.0000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 781.8500 1119.4800 781.9500 1120.0000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 777.8500 1119.4800 777.9500 1120.0000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 773.8500 1119.4800 773.9500 1120.0000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 769.8500 1119.4800 769.9500 1120.0000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 765.8500 1119.4800 765.9500 1120.0000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 761.8500 1119.4800 761.9500 1120.0000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 757.8500 1119.4800 757.9500 1120.0000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 753.8500 1119.4800 753.9500 1120.0000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 749.8500 1119.4800 749.9500 1120.0000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 745.8500 1119.4800 745.9500 1120.0000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 741.8500 1119.4800 741.9500 1120.0000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 737.8500 1119.4800 737.9500 1120.0000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 733.8500 1119.4800 733.9500 1120.0000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 729.8500 1119.4800 729.9500 1120.0000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 725.8500 1119.4800 725.9500 1120.0000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 721.8500 1119.4800 721.9500 1120.0000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 717.8500 1119.4800 717.9500 1120.0000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 713.8500 1119.4800 713.9500 1120.0000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 709.8500 1119.4800 709.9500 1120.0000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 705.8500 1119.4800 705.9500 1120.0000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 701.8500 1119.4800 701.9500 1120.0000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 697.8500 1119.4800 697.9500 1120.0000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 693.8500 1119.4800 693.9500 1120.0000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 689.8500 1119.4800 689.9500 1120.0000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 685.8500 1119.4800 685.9500 1120.0000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 681.8500 1119.4800 681.9500 1120.0000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 677.8500 1119.4800 677.9500 1120.0000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 673.8500 1119.4800 673.9500 1120.0000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 669.8500 1119.4800 669.9500 1120.0000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.8500 1119.4800 665.9500 1120.0000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 661.8500 1119.4800 661.9500 1120.0000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 657.8500 1119.4800 657.9500 1120.0000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 653.8500 1119.4800 653.9500 1120.0000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 649.8500 1119.4800 649.9500 1120.0000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 645.8500 1119.4800 645.9500 1120.0000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 641.8500 1119.4800 641.9500 1120.0000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 637.8500 1119.4800 637.9500 1120.0000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 633.8500 1119.4800 633.9500 1120.0000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 629.8500 1119.4800 629.9500 1120.0000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 625.8500 1119.4800 625.9500 1120.0000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 621.8500 1119.4800 621.9500 1120.0000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 617.8500 1119.4800 617.9500 1120.0000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 613.8500 1119.4800 613.9500 1120.0000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 609.8500 1119.4800 609.9500 1120.0000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 605.8500 1119.4800 605.9500 1120.0000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 601.8500 1119.4800 601.9500 1120.0000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 597.8500 1119.4800 597.9500 1120.0000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 593.8500 1119.4800 593.9500 1120.0000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 589.8500 1119.4800 589.9500 1120.0000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 585.8500 1119.4800 585.9500 1120.0000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 581.8500 1119.4800 581.9500 1120.0000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 577.8500 1119.4800 577.9500 1120.0000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 573.8500 1119.4800 573.9500 1120.0000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 569.8500 1119.4800 569.9500 1120.0000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 565.8500 1119.4800 565.9500 1120.0000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 561.8500 1119.4800 561.9500 1120.0000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 557.8500 1119.4800 557.9500 1120.0000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 553.8500 1119.4800 553.9500 1120.0000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 549.8500 1119.4800 549.9500 1120.0000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 545.8500 1119.4800 545.9500 1120.0000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 541.8500 1119.4800 541.9500 1120.0000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 537.8500 1119.4800 537.9500 1120.0000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 533.8500 1119.4800 533.9500 1120.0000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 529.8500 1119.4800 529.9500 1120.0000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 525.8500 1119.4800 525.9500 1120.0000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 521.8500 1119.4800 521.9500 1120.0000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 517.8500 1119.4800 517.9500 1120.0000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 513.8500 1119.4800 513.9500 1120.0000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 509.8500 1119.4800 509.9500 1120.0000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 505.8500 1119.4800 505.9500 1120.0000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 501.8500 1119.4800 501.9500 1120.0000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 497.8500 1119.4800 497.9500 1120.0000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 493.8500 1119.4800 493.9500 1120.0000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 489.8500 1119.4800 489.9500 1120.0000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 485.8500 1119.4800 485.9500 1120.0000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 481.8500 1119.4800 481.9500 1120.0000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 477.8500 1119.4800 477.9500 1120.0000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 473.8500 1119.4800 473.9500 1120.0000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 469.8500 1119.4800 469.9500 1120.0000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 465.8500 1119.4800 465.9500 1120.0000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 461.8500 1119.4800 461.9500 1120.0000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.8500 1119.4800 457.9500 1120.0000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 453.8500 1119.4800 453.9500 1120.0000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.8500 1119.4800 449.9500 1120.0000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.8500 1119.4800 445.9500 1120.0000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.8500 1119.4800 441.9500 1120.0000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 437.8500 1119.4800 437.9500 1120.0000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.8500 1119.4800 433.9500 1120.0000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 429.8500 1119.4800 429.9500 1120.0000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.8500 1119.4800 425.9500 1120.0000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 421.8500 1119.4800 421.9500 1120.0000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.8500 1119.4800 417.9500 1120.0000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 413.8500 1119.4800 413.9500 1120.0000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 409.8500 1119.4800 409.9500 1120.0000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.8500 1119.4800 405.9500 1120.0000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 401.8500 1119.4800 401.9500 1120.0000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.8500 1119.4800 397.9500 1120.0000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 393.8500 1119.4800 393.9500 1120.0000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.8500 1119.4800 389.9500 1120.0000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.8500 1119.4800 385.9500 1120.0000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.8500 1119.4800 381.9500 1120.0000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 377.8500 1119.4800 377.9500 1120.0000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.8500 1119.4800 373.9500 1120.0000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.8500 1119.4800 369.9500 1120.0000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.8500 1119.4800 365.9500 1120.0000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.8500 1119.4800 361.9500 1120.0000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.8500 1119.4800 357.9500 1120.0000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.8500 1119.4800 353.9500 1120.0000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.8500 1119.4800 349.9500 1120.0000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.8500 1119.4800 345.9500 1120.0000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.8500 1119.4800 341.9500 1120.0000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.8500 1119.4800 337.9500 1120.0000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.8500 1119.4800 333.9500 1120.0000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.8500 1119.4800 329.9500 1120.0000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.8500 1119.4800 325.9500 1120.0000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.8500 1119.4800 321.9500 1120.0000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.8500 1119.4800 317.9500 1120.0000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.8500 1119.4800 313.9500 1120.0000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.8500 1119.4800 309.9500 1120.0000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.8500 1119.4800 305.9500 1120.0000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 301.8500 1119.4800 301.9500 1120.0000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.8500 1119.4800 297.9500 1120.0000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 293.8500 1119.4800 293.9500 1120.0000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.8500 1119.4800 289.9500 1120.0000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.8500 1119.4800 285.9500 1120.0000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.8500 1119.4800 281.9500 1120.0000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.8500 1119.4800 277.9500 1120.0000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.8500 1119.4800 273.9500 1120.0000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 269.8500 1119.4800 269.9500 1120.0000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.8500 1119.4800 265.9500 1120.0000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.8500 1119.4800 261.9500 1120.0000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 257.8500 1119.4800 257.9500 1120.0000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 253.8500 1119.4800 253.9500 1120.0000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 249.8500 1119.4800 249.9500 1120.0000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.8500 1119.4800 245.9500 1120.0000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.8500 1119.4800 241.9500 1120.0000 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 587.7500 0.5200 587.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 583.7500 0.5200 583.8500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 579.7500 0.5200 579.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 575.7500 0.5200 575.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 571.7500 0.5200 571.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 567.7500 0.5200 567.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 563.7500 0.5200 563.8500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 559.7500 0.5200 559.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 555.7500 0.5200 555.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 551.7500 0.5200 551.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 547.7500 0.5200 547.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 543.7500 0.5200 543.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 539.7500 0.5200 539.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 535.7500 0.5200 535.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 531.7500 0.5200 531.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 527.7500 0.5200 527.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 523.7500 0.5200 523.8500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 595.7500 0.5200 595.8500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1120.0000 1120.0000 ;
    LAYER M2 ;
      RECT 878.0500 1119.3800 1120.0000 1120.0000 ;
      RECT 874.0500 1119.3800 877.7500 1120.0000 ;
      RECT 870.0500 1119.3800 873.7500 1120.0000 ;
      RECT 866.0500 1119.3800 869.7500 1120.0000 ;
      RECT 862.0500 1119.3800 865.7500 1120.0000 ;
      RECT 858.0500 1119.3800 861.7500 1120.0000 ;
      RECT 854.0500 1119.3800 857.7500 1120.0000 ;
      RECT 850.0500 1119.3800 853.7500 1120.0000 ;
      RECT 846.0500 1119.3800 849.7500 1120.0000 ;
      RECT 842.0500 1119.3800 845.7500 1120.0000 ;
      RECT 838.0500 1119.3800 841.7500 1120.0000 ;
      RECT 834.0500 1119.3800 837.7500 1120.0000 ;
      RECT 830.0500 1119.3800 833.7500 1120.0000 ;
      RECT 826.0500 1119.3800 829.7500 1120.0000 ;
      RECT 822.0500 1119.3800 825.7500 1120.0000 ;
      RECT 818.0500 1119.3800 821.7500 1120.0000 ;
      RECT 814.0500 1119.3800 817.7500 1120.0000 ;
      RECT 810.0500 1119.3800 813.7500 1120.0000 ;
      RECT 806.0500 1119.3800 809.7500 1120.0000 ;
      RECT 802.0500 1119.3800 805.7500 1120.0000 ;
      RECT 798.0500 1119.3800 801.7500 1120.0000 ;
      RECT 794.0500 1119.3800 797.7500 1120.0000 ;
      RECT 790.0500 1119.3800 793.7500 1120.0000 ;
      RECT 786.0500 1119.3800 789.7500 1120.0000 ;
      RECT 782.0500 1119.3800 785.7500 1120.0000 ;
      RECT 778.0500 1119.3800 781.7500 1120.0000 ;
      RECT 774.0500 1119.3800 777.7500 1120.0000 ;
      RECT 770.0500 1119.3800 773.7500 1120.0000 ;
      RECT 766.0500 1119.3800 769.7500 1120.0000 ;
      RECT 762.0500 1119.3800 765.7500 1120.0000 ;
      RECT 758.0500 1119.3800 761.7500 1120.0000 ;
      RECT 754.0500 1119.3800 757.7500 1120.0000 ;
      RECT 750.0500 1119.3800 753.7500 1120.0000 ;
      RECT 746.0500 1119.3800 749.7500 1120.0000 ;
      RECT 742.0500 1119.3800 745.7500 1120.0000 ;
      RECT 738.0500 1119.3800 741.7500 1120.0000 ;
      RECT 734.0500 1119.3800 737.7500 1120.0000 ;
      RECT 730.0500 1119.3800 733.7500 1120.0000 ;
      RECT 726.0500 1119.3800 729.7500 1120.0000 ;
      RECT 722.0500 1119.3800 725.7500 1120.0000 ;
      RECT 718.0500 1119.3800 721.7500 1120.0000 ;
      RECT 714.0500 1119.3800 717.7500 1120.0000 ;
      RECT 710.0500 1119.3800 713.7500 1120.0000 ;
      RECT 706.0500 1119.3800 709.7500 1120.0000 ;
      RECT 702.0500 1119.3800 705.7500 1120.0000 ;
      RECT 698.0500 1119.3800 701.7500 1120.0000 ;
      RECT 694.0500 1119.3800 697.7500 1120.0000 ;
      RECT 690.0500 1119.3800 693.7500 1120.0000 ;
      RECT 686.0500 1119.3800 689.7500 1120.0000 ;
      RECT 682.0500 1119.3800 685.7500 1120.0000 ;
      RECT 678.0500 1119.3800 681.7500 1120.0000 ;
      RECT 674.0500 1119.3800 677.7500 1120.0000 ;
      RECT 670.0500 1119.3800 673.7500 1120.0000 ;
      RECT 666.0500 1119.3800 669.7500 1120.0000 ;
      RECT 662.0500 1119.3800 665.7500 1120.0000 ;
      RECT 658.0500 1119.3800 661.7500 1120.0000 ;
      RECT 654.0500 1119.3800 657.7500 1120.0000 ;
      RECT 650.0500 1119.3800 653.7500 1120.0000 ;
      RECT 646.0500 1119.3800 649.7500 1120.0000 ;
      RECT 642.0500 1119.3800 645.7500 1120.0000 ;
      RECT 638.0500 1119.3800 641.7500 1120.0000 ;
      RECT 634.0500 1119.3800 637.7500 1120.0000 ;
      RECT 630.0500 1119.3800 633.7500 1120.0000 ;
      RECT 626.0500 1119.3800 629.7500 1120.0000 ;
      RECT 622.0500 1119.3800 625.7500 1120.0000 ;
      RECT 618.0500 1119.3800 621.7500 1120.0000 ;
      RECT 614.0500 1119.3800 617.7500 1120.0000 ;
      RECT 610.0500 1119.3800 613.7500 1120.0000 ;
      RECT 606.0500 1119.3800 609.7500 1120.0000 ;
      RECT 602.0500 1119.3800 605.7500 1120.0000 ;
      RECT 598.0500 1119.3800 601.7500 1120.0000 ;
      RECT 594.0500 1119.3800 597.7500 1120.0000 ;
      RECT 590.0500 1119.3800 593.7500 1120.0000 ;
      RECT 586.0500 1119.3800 589.7500 1120.0000 ;
      RECT 582.0500 1119.3800 585.7500 1120.0000 ;
      RECT 578.0500 1119.3800 581.7500 1120.0000 ;
      RECT 574.0500 1119.3800 577.7500 1120.0000 ;
      RECT 570.0500 1119.3800 573.7500 1120.0000 ;
      RECT 566.0500 1119.3800 569.7500 1120.0000 ;
      RECT 562.0500 1119.3800 565.7500 1120.0000 ;
      RECT 558.0500 1119.3800 561.7500 1120.0000 ;
      RECT 554.0500 1119.3800 557.7500 1120.0000 ;
      RECT 550.0500 1119.3800 553.7500 1120.0000 ;
      RECT 546.0500 1119.3800 549.7500 1120.0000 ;
      RECT 542.0500 1119.3800 545.7500 1120.0000 ;
      RECT 538.0500 1119.3800 541.7500 1120.0000 ;
      RECT 534.0500 1119.3800 537.7500 1120.0000 ;
      RECT 530.0500 1119.3800 533.7500 1120.0000 ;
      RECT 526.0500 1119.3800 529.7500 1120.0000 ;
      RECT 522.0500 1119.3800 525.7500 1120.0000 ;
      RECT 518.0500 1119.3800 521.7500 1120.0000 ;
      RECT 514.0500 1119.3800 517.7500 1120.0000 ;
      RECT 510.0500 1119.3800 513.7500 1120.0000 ;
      RECT 506.0500 1119.3800 509.7500 1120.0000 ;
      RECT 502.0500 1119.3800 505.7500 1120.0000 ;
      RECT 498.0500 1119.3800 501.7500 1120.0000 ;
      RECT 494.0500 1119.3800 497.7500 1120.0000 ;
      RECT 490.0500 1119.3800 493.7500 1120.0000 ;
      RECT 486.0500 1119.3800 489.7500 1120.0000 ;
      RECT 482.0500 1119.3800 485.7500 1120.0000 ;
      RECT 478.0500 1119.3800 481.7500 1120.0000 ;
      RECT 474.0500 1119.3800 477.7500 1120.0000 ;
      RECT 470.0500 1119.3800 473.7500 1120.0000 ;
      RECT 466.0500 1119.3800 469.7500 1120.0000 ;
      RECT 462.0500 1119.3800 465.7500 1120.0000 ;
      RECT 458.0500 1119.3800 461.7500 1120.0000 ;
      RECT 454.0500 1119.3800 457.7500 1120.0000 ;
      RECT 450.0500 1119.3800 453.7500 1120.0000 ;
      RECT 446.0500 1119.3800 449.7500 1120.0000 ;
      RECT 442.0500 1119.3800 445.7500 1120.0000 ;
      RECT 438.0500 1119.3800 441.7500 1120.0000 ;
      RECT 434.0500 1119.3800 437.7500 1120.0000 ;
      RECT 430.0500 1119.3800 433.7500 1120.0000 ;
      RECT 426.0500 1119.3800 429.7500 1120.0000 ;
      RECT 422.0500 1119.3800 425.7500 1120.0000 ;
      RECT 418.0500 1119.3800 421.7500 1120.0000 ;
      RECT 414.0500 1119.3800 417.7500 1120.0000 ;
      RECT 410.0500 1119.3800 413.7500 1120.0000 ;
      RECT 406.0500 1119.3800 409.7500 1120.0000 ;
      RECT 402.0500 1119.3800 405.7500 1120.0000 ;
      RECT 398.0500 1119.3800 401.7500 1120.0000 ;
      RECT 394.0500 1119.3800 397.7500 1120.0000 ;
      RECT 390.0500 1119.3800 393.7500 1120.0000 ;
      RECT 386.0500 1119.3800 389.7500 1120.0000 ;
      RECT 382.0500 1119.3800 385.7500 1120.0000 ;
      RECT 378.0500 1119.3800 381.7500 1120.0000 ;
      RECT 374.0500 1119.3800 377.7500 1120.0000 ;
      RECT 370.0500 1119.3800 373.7500 1120.0000 ;
      RECT 366.0500 1119.3800 369.7500 1120.0000 ;
      RECT 362.0500 1119.3800 365.7500 1120.0000 ;
      RECT 358.0500 1119.3800 361.7500 1120.0000 ;
      RECT 354.0500 1119.3800 357.7500 1120.0000 ;
      RECT 350.0500 1119.3800 353.7500 1120.0000 ;
      RECT 346.0500 1119.3800 349.7500 1120.0000 ;
      RECT 342.0500 1119.3800 345.7500 1120.0000 ;
      RECT 338.0500 1119.3800 341.7500 1120.0000 ;
      RECT 334.0500 1119.3800 337.7500 1120.0000 ;
      RECT 330.0500 1119.3800 333.7500 1120.0000 ;
      RECT 326.0500 1119.3800 329.7500 1120.0000 ;
      RECT 322.0500 1119.3800 325.7500 1120.0000 ;
      RECT 318.0500 1119.3800 321.7500 1120.0000 ;
      RECT 314.0500 1119.3800 317.7500 1120.0000 ;
      RECT 310.0500 1119.3800 313.7500 1120.0000 ;
      RECT 306.0500 1119.3800 309.7500 1120.0000 ;
      RECT 302.0500 1119.3800 305.7500 1120.0000 ;
      RECT 298.0500 1119.3800 301.7500 1120.0000 ;
      RECT 294.0500 1119.3800 297.7500 1120.0000 ;
      RECT 290.0500 1119.3800 293.7500 1120.0000 ;
      RECT 286.0500 1119.3800 289.7500 1120.0000 ;
      RECT 282.0500 1119.3800 285.7500 1120.0000 ;
      RECT 278.0500 1119.3800 281.7500 1120.0000 ;
      RECT 274.0500 1119.3800 277.7500 1120.0000 ;
      RECT 270.0500 1119.3800 273.7500 1120.0000 ;
      RECT 266.0500 1119.3800 269.7500 1120.0000 ;
      RECT 262.0500 1119.3800 265.7500 1120.0000 ;
      RECT 258.0500 1119.3800 261.7500 1120.0000 ;
      RECT 254.0500 1119.3800 257.7500 1120.0000 ;
      RECT 250.0500 1119.3800 253.7500 1120.0000 ;
      RECT 246.0500 1119.3800 249.7500 1120.0000 ;
      RECT 242.0500 1119.3800 245.7500 1120.0000 ;
      RECT 0.0000 1119.3800 241.7500 1120.0000 ;
      RECT 0.0000 0.6200 1120.0000 1119.3800 ;
      RECT 686.0500 0.0000 1120.0000 0.6200 ;
      RECT 682.0500 0.0000 685.7500 0.6200 ;
      RECT 678.0500 0.0000 681.7500 0.6200 ;
      RECT 674.0500 0.0000 677.7500 0.6200 ;
      RECT 670.0500 0.0000 673.7500 0.6200 ;
      RECT 666.0500 0.0000 669.7500 0.6200 ;
      RECT 662.0500 0.0000 665.7500 0.6200 ;
      RECT 658.0500 0.0000 661.7500 0.6200 ;
      RECT 654.0500 0.0000 657.7500 0.6200 ;
      RECT 650.0500 0.0000 653.7500 0.6200 ;
      RECT 646.0500 0.0000 649.7500 0.6200 ;
      RECT 642.0500 0.0000 645.7500 0.6200 ;
      RECT 638.0500 0.0000 641.7500 0.6200 ;
      RECT 634.0500 0.0000 637.7500 0.6200 ;
      RECT 630.0500 0.0000 633.7500 0.6200 ;
      RECT 626.0500 0.0000 629.7500 0.6200 ;
      RECT 622.0500 0.0000 625.7500 0.6200 ;
      RECT 618.0500 0.0000 621.7500 0.6200 ;
      RECT 614.0500 0.0000 617.7500 0.6200 ;
      RECT 610.0500 0.0000 613.7500 0.6200 ;
      RECT 606.0500 0.0000 609.7500 0.6200 ;
      RECT 602.0500 0.0000 605.7500 0.6200 ;
      RECT 598.0500 0.0000 601.7500 0.6200 ;
      RECT 594.0500 0.0000 597.7500 0.6200 ;
      RECT 590.0500 0.0000 593.7500 0.6200 ;
      RECT 586.0500 0.0000 589.7500 0.6200 ;
      RECT 582.0500 0.0000 585.7500 0.6200 ;
      RECT 578.0500 0.0000 581.7500 0.6200 ;
      RECT 574.0500 0.0000 577.7500 0.6200 ;
      RECT 570.0500 0.0000 573.7500 0.6200 ;
      RECT 566.0500 0.0000 569.7500 0.6200 ;
      RECT 562.0500 0.0000 565.7500 0.6200 ;
      RECT 558.0500 0.0000 561.7500 0.6200 ;
      RECT 554.0500 0.0000 557.7500 0.6200 ;
      RECT 550.0500 0.0000 553.7500 0.6200 ;
      RECT 546.0500 0.0000 549.7500 0.6200 ;
      RECT 542.0500 0.0000 545.7500 0.6200 ;
      RECT 538.0500 0.0000 541.7500 0.6200 ;
      RECT 534.0500 0.0000 537.7500 0.6200 ;
      RECT 530.0500 0.0000 533.7500 0.6200 ;
      RECT 526.0500 0.0000 529.7500 0.6200 ;
      RECT 522.0500 0.0000 525.7500 0.6200 ;
      RECT 518.0500 0.0000 521.7500 0.6200 ;
      RECT 514.0500 0.0000 517.7500 0.6200 ;
      RECT 510.0500 0.0000 513.7500 0.6200 ;
      RECT 506.0500 0.0000 509.7500 0.6200 ;
      RECT 502.0500 0.0000 505.7500 0.6200 ;
      RECT 498.0500 0.0000 501.7500 0.6200 ;
      RECT 494.0500 0.0000 497.7500 0.6200 ;
      RECT 490.0500 0.0000 493.7500 0.6200 ;
      RECT 486.0500 0.0000 489.7500 0.6200 ;
      RECT 482.0500 0.0000 485.7500 0.6200 ;
      RECT 478.0500 0.0000 481.7500 0.6200 ;
      RECT 474.0500 0.0000 477.7500 0.6200 ;
      RECT 470.0500 0.0000 473.7500 0.6200 ;
      RECT 466.0500 0.0000 469.7500 0.6200 ;
      RECT 462.0500 0.0000 465.7500 0.6200 ;
      RECT 458.0500 0.0000 461.7500 0.6200 ;
      RECT 454.0500 0.0000 457.7500 0.6200 ;
      RECT 450.0500 0.0000 453.7500 0.6200 ;
      RECT 446.0500 0.0000 449.7500 0.6200 ;
      RECT 442.0500 0.0000 445.7500 0.6200 ;
      RECT 438.0500 0.0000 441.7500 0.6200 ;
      RECT 434.0500 0.0000 437.7500 0.6200 ;
      RECT 0.0000 0.0000 433.7500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 595.9500 1120.0000 1120.0000 ;
      RECT 0.6200 595.6500 1120.0000 595.9500 ;
      RECT 0.0000 591.9500 1120.0000 595.6500 ;
      RECT 0.6200 591.6500 1120.0000 591.9500 ;
      RECT 0.0000 587.9500 1120.0000 591.6500 ;
      RECT 0.6200 587.6500 1120.0000 587.9500 ;
      RECT 0.0000 583.9500 1120.0000 587.6500 ;
      RECT 0.6200 583.6500 1120.0000 583.9500 ;
      RECT 0.0000 579.9500 1120.0000 583.6500 ;
      RECT 0.6200 579.6500 1120.0000 579.9500 ;
      RECT 0.0000 575.9500 1120.0000 579.6500 ;
      RECT 0.6200 575.6500 1120.0000 575.9500 ;
      RECT 0.0000 571.9500 1120.0000 575.6500 ;
      RECT 0.6200 571.6500 1120.0000 571.9500 ;
      RECT 0.0000 567.9500 1120.0000 571.6500 ;
      RECT 0.6200 567.6500 1120.0000 567.9500 ;
      RECT 0.0000 563.9500 1120.0000 567.6500 ;
      RECT 0.6200 563.6500 1120.0000 563.9500 ;
      RECT 0.0000 559.9500 1120.0000 563.6500 ;
      RECT 0.6200 559.6500 1120.0000 559.9500 ;
      RECT 0.0000 555.9500 1120.0000 559.6500 ;
      RECT 0.6200 555.6500 1120.0000 555.9500 ;
      RECT 0.0000 551.9500 1120.0000 555.6500 ;
      RECT 0.6200 551.6500 1120.0000 551.9500 ;
      RECT 0.0000 547.9500 1120.0000 551.6500 ;
      RECT 0.6200 547.6500 1120.0000 547.9500 ;
      RECT 0.0000 543.9500 1120.0000 547.6500 ;
      RECT 0.6200 543.6500 1120.0000 543.9500 ;
      RECT 0.0000 539.9500 1120.0000 543.6500 ;
      RECT 0.6200 539.6500 1120.0000 539.9500 ;
      RECT 0.0000 535.9500 1120.0000 539.6500 ;
      RECT 0.6200 535.6500 1120.0000 535.9500 ;
      RECT 0.0000 531.9500 1120.0000 535.6500 ;
      RECT 0.6200 531.6500 1120.0000 531.9500 ;
      RECT 0.0000 527.9500 1120.0000 531.6500 ;
      RECT 0.6200 527.6500 1120.0000 527.9500 ;
      RECT 0.0000 523.9500 1120.0000 527.6500 ;
      RECT 0.6200 523.6500 1120.0000 523.9500 ;
      RECT 0.0000 0.0000 1120.0000 523.6500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 1120.0000 1120.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 1120.0000 1120.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 1120.0000 1120.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 1120.0000 1120.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 1120.0000 1120.0000 ;
  END
END core

END LIBRARY
