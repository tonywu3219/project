##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 20:00:54 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 1220.0000 BY 1220.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 567.7500 0.5200 567.8500 ;
    END
  END clk
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.8500 1219.4800 287.9500 1220.0000 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.8500 1219.4800 283.9500 1220.0000 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.8500 1219.4800 279.9500 1220.0000 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.8500 1219.4800 275.9500 1220.0000 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.8500 1219.4800 271.9500 1220.0000 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.8500 1219.4800 267.9500 1220.0000 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.8500 1219.4800 263.9500 1220.0000 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.8500 1219.4800 259.9500 1220.0000 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.8500 1219.4800 255.9500 1220.0000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.8500 1219.4800 251.9500 1220.0000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.8500 1219.4800 247.9500 1220.0000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.8500 1219.4800 243.9500 1220.0000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 239.8500 1219.4800 239.9500 1220.0000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.8500 1219.4800 235.9500 1220.0000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.8500 1219.4800 231.9500 1220.0000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.8500 1219.4800 227.9500 1220.0000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.8500 1219.4800 223.9500 1220.0000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.8500 1219.4800 219.9500 1220.0000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.8500 1219.4800 215.9500 1220.0000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.8500 1219.4800 211.9500 1220.0000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.8500 1219.4800 207.9500 1220.0000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.8500 1219.4800 203.9500 1220.0000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.8500 1219.4800 199.9500 1220.0000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.8500 1219.4800 195.9500 1220.0000 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 735.8500 0.0000 735.9500 0.5200 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 731.8500 0.0000 731.9500 0.5200 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 727.8500 0.0000 727.9500 0.5200 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 723.8500 0.0000 723.9500 0.5200 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 719.8500 0.0000 719.9500 0.5200 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 715.8500 0.0000 715.9500 0.5200 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 711.8500 0.0000 711.9500 0.5200 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 707.8500 0.0000 707.9500 0.5200 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 703.8500 0.0000 703.9500 0.5200 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 699.8500 0.0000 699.9500 0.5200 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 695.8500 0.0000 695.9500 0.5200 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 691.8500 0.0000 691.9500 0.5200 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 687.8500 0.0000 687.9500 0.5200 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 683.8500 0.0000 683.9500 0.5200 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 679.8500 0.0000 679.9500 0.5200 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 675.8500 0.0000 675.9500 0.5200 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 671.8500 0.0000 671.9500 0.5200 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 667.8500 0.0000 667.9500 0.5200 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 663.8500 0.0000 663.9500 0.5200 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 659.8500 0.0000 659.9500 0.5200 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 655.8500 0.0000 655.9500 0.5200 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 651.8500 0.0000 651.9500 0.5200 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 647.8500 0.0000 647.9500 0.5200 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 643.8500 0.0000 643.9500 0.5200 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 639.8500 0.0000 639.9500 0.5200 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 635.8500 0.0000 635.9500 0.5200 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 631.8500 0.0000 631.9500 0.5200 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 627.8500 0.0000 627.9500 0.5200 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 623.8500 0.0000 623.9500 0.5200 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 619.8500 0.0000 619.9500 0.5200 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 615.8500 0.0000 615.9500 0.5200 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 611.8500 0.0000 611.9500 0.5200 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 607.8500 0.0000 607.9500 0.5200 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 603.8500 0.0000 603.9500 0.5200 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 599.8500 0.0000 599.9500 0.5200 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 595.8500 0.0000 595.9500 0.5200 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 591.8500 0.0000 591.9500 0.5200 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 587.8500 0.0000 587.9500 0.5200 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 583.8500 0.0000 583.9500 0.5200 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 579.8500 0.0000 579.9500 0.5200 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 575.8500 0.0000 575.9500 0.5200 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 571.8500 0.0000 571.9500 0.5200 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 567.8500 0.0000 567.9500 0.5200 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 563.8500 0.0000 563.9500 0.5200 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 559.8500 0.0000 559.9500 0.5200 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 555.8500 0.0000 555.9500 0.5200 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 551.8500 0.0000 551.9500 0.5200 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 547.8500 0.0000 547.9500 0.5200 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 543.8500 0.0000 543.9500 0.5200 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 539.8500 0.0000 539.9500 0.5200 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 535.8500 0.0000 535.9500 0.5200 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 531.8500 0.0000 531.9500 0.5200 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 527.8500 0.0000 527.9500 0.5200 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 523.8500 0.0000 523.9500 0.5200 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 519.8500 0.0000 519.9500 0.5200 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 515.8500 0.0000 515.9500 0.5200 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 511.8500 0.0000 511.9500 0.5200 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.8500 0.0000 507.9500 0.5200 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 503.8500 0.0000 503.9500 0.5200 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 499.8500 0.0000 499.9500 0.5200 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 495.8500 0.0000 495.9500 0.5200 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 491.8500 0.0000 491.9500 0.5200 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 487.8500 0.0000 487.9500 0.5200 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 483.8500 0.0000 483.9500 0.5200 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1023.8500 1219.4800 1023.9500 1220.0000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1019.8500 1219.4800 1019.9500 1220.0000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1015.8500 1219.4800 1015.9500 1220.0000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1011.8500 1219.4800 1011.9500 1220.0000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1007.8500 1219.4800 1007.9500 1220.0000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1003.8500 1219.4800 1003.9500 1220.0000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 999.8500 1219.4800 999.9500 1220.0000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 995.8500 1219.4800 995.9500 1220.0000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 991.8500 1219.4800 991.9500 1220.0000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 987.8500 1219.4800 987.9500 1220.0000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 983.8500 1219.4800 983.9500 1220.0000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 979.8500 1219.4800 979.9500 1220.0000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 975.8500 1219.4800 975.9500 1220.0000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 971.8500 1219.4800 971.9500 1220.0000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 967.8500 1219.4800 967.9500 1220.0000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 963.8500 1219.4800 963.9500 1220.0000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 959.8500 1219.4800 959.9500 1220.0000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 955.8500 1219.4800 955.9500 1220.0000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 951.8500 1219.4800 951.9500 1220.0000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 947.8500 1219.4800 947.9500 1220.0000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 943.8500 1219.4800 943.9500 1220.0000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 939.8500 1219.4800 939.9500 1220.0000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 935.8500 1219.4800 935.9500 1220.0000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 931.8500 1219.4800 931.9500 1220.0000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 927.8500 1219.4800 927.9500 1220.0000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 923.8500 1219.4800 923.9500 1220.0000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 919.8500 1219.4800 919.9500 1220.0000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 915.8500 1219.4800 915.9500 1220.0000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 911.8500 1219.4800 911.9500 1220.0000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 907.8500 1219.4800 907.9500 1220.0000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 903.8500 1219.4800 903.9500 1220.0000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 899.8500 1219.4800 899.9500 1220.0000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 895.8500 1219.4800 895.9500 1220.0000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 891.8500 1219.4800 891.9500 1220.0000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 887.8500 1219.4800 887.9500 1220.0000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 883.8500 1219.4800 883.9500 1220.0000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 879.8500 1219.4800 879.9500 1220.0000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 875.8500 1219.4800 875.9500 1220.0000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 871.8500 1219.4800 871.9500 1220.0000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 867.8500 1219.4800 867.9500 1220.0000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 863.8500 1219.4800 863.9500 1220.0000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 859.8500 1219.4800 859.9500 1220.0000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 855.8500 1219.4800 855.9500 1220.0000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 851.8500 1219.4800 851.9500 1220.0000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 847.8500 1219.4800 847.9500 1220.0000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 843.8500 1219.4800 843.9500 1220.0000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 839.8500 1219.4800 839.9500 1220.0000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 835.8500 1219.4800 835.9500 1220.0000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 831.8500 1219.4800 831.9500 1220.0000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 827.8500 1219.4800 827.9500 1220.0000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 823.8500 1219.4800 823.9500 1220.0000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 819.8500 1219.4800 819.9500 1220.0000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 815.8500 1219.4800 815.9500 1220.0000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 811.8500 1219.4800 811.9500 1220.0000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 807.8500 1219.4800 807.9500 1220.0000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 803.8500 1219.4800 803.9500 1220.0000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 799.8500 1219.4800 799.9500 1220.0000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 795.8500 1219.4800 795.9500 1220.0000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 791.8500 1219.4800 791.9500 1220.0000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 787.8500 1219.4800 787.9500 1220.0000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 783.8500 1219.4800 783.9500 1220.0000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 779.8500 1219.4800 779.9500 1220.0000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 775.8500 1219.4800 775.9500 1220.0000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 771.8500 1219.4800 771.9500 1220.0000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 767.8500 1219.4800 767.9500 1220.0000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 763.8500 1219.4800 763.9500 1220.0000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 759.8500 1219.4800 759.9500 1220.0000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 755.8500 1219.4800 755.9500 1220.0000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 751.8500 1219.4800 751.9500 1220.0000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 747.8500 1219.4800 747.9500 1220.0000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 743.8500 1219.4800 743.9500 1220.0000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 739.8500 1219.4800 739.9500 1220.0000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 735.8500 1219.4800 735.9500 1220.0000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 731.8500 1219.4800 731.9500 1220.0000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 727.8500 1219.4800 727.9500 1220.0000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 723.8500 1219.4800 723.9500 1220.0000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 719.8500 1219.4800 719.9500 1220.0000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 715.8500 1219.4800 715.9500 1220.0000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 711.8500 1219.4800 711.9500 1220.0000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 707.8500 1219.4800 707.9500 1220.0000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 703.8500 1219.4800 703.9500 1220.0000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 699.8500 1219.4800 699.9500 1220.0000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 695.8500 1219.4800 695.9500 1220.0000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 691.8500 1219.4800 691.9500 1220.0000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 687.8500 1219.4800 687.9500 1220.0000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 683.8500 1219.4800 683.9500 1220.0000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 679.8500 1219.4800 679.9500 1220.0000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 675.8500 1219.4800 675.9500 1220.0000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 671.8500 1219.4800 671.9500 1220.0000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 667.8500 1219.4800 667.9500 1220.0000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 663.8500 1219.4800 663.9500 1220.0000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 659.8500 1219.4800 659.9500 1220.0000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 655.8500 1219.4800 655.9500 1220.0000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 651.8500 1219.4800 651.9500 1220.0000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 647.8500 1219.4800 647.9500 1220.0000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 643.8500 1219.4800 643.9500 1220.0000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 639.8500 1219.4800 639.9500 1220.0000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 635.8500 1219.4800 635.9500 1220.0000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 631.8500 1219.4800 631.9500 1220.0000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 627.8500 1219.4800 627.9500 1220.0000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 623.8500 1219.4800 623.9500 1220.0000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 619.8500 1219.4800 619.9500 1220.0000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 615.8500 1219.4800 615.9500 1220.0000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 611.8500 1219.4800 611.9500 1220.0000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 607.8500 1219.4800 607.9500 1220.0000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 603.8500 1219.4800 603.9500 1220.0000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 599.8500 1219.4800 599.9500 1220.0000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 595.8500 1219.4800 595.9500 1220.0000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 591.8500 1219.4800 591.9500 1220.0000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 587.8500 1219.4800 587.9500 1220.0000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 583.8500 1219.4800 583.9500 1220.0000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 579.8500 1219.4800 579.9500 1220.0000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 575.8500 1219.4800 575.9500 1220.0000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 571.8500 1219.4800 571.9500 1220.0000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 567.8500 1219.4800 567.9500 1220.0000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 563.8500 1219.4800 563.9500 1220.0000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 559.8500 1219.4800 559.9500 1220.0000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 555.8500 1219.4800 555.9500 1220.0000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 551.8500 1219.4800 551.9500 1220.0000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 547.8500 1219.4800 547.9500 1220.0000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 543.8500 1219.4800 543.9500 1220.0000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 539.8500 1219.4800 539.9500 1220.0000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 535.8500 1219.4800 535.9500 1220.0000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 531.8500 1219.4800 531.9500 1220.0000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 527.8500 1219.4800 527.9500 1220.0000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 523.8500 1219.4800 523.9500 1220.0000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 519.8500 1219.4800 519.9500 1220.0000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 515.8500 1219.4800 515.9500 1220.0000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 511.8500 1219.4800 511.9500 1220.0000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.8500 1219.4800 507.9500 1220.0000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 503.8500 1219.4800 503.9500 1220.0000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 499.8500 1219.4800 499.9500 1220.0000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 495.8500 1219.4800 495.9500 1220.0000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 491.8500 1219.4800 491.9500 1220.0000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 487.8500 1219.4800 487.9500 1220.0000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 483.8500 1219.4800 483.9500 1220.0000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 479.8500 1219.4800 479.9500 1220.0000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 475.8500 1219.4800 475.9500 1220.0000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 471.8500 1219.4800 471.9500 1220.0000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 467.8500 1219.4800 467.9500 1220.0000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.8500 1219.4800 463.9500 1220.0000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 459.8500 1219.4800 459.9500 1220.0000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.8500 1219.4800 455.9500 1220.0000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.8500 1219.4800 451.9500 1220.0000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.8500 1219.4800 447.9500 1220.0000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.8500 1219.4800 443.9500 1220.0000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.8500 1219.4800 439.9500 1220.0000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.8500 1219.4800 435.9500 1220.0000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.8500 1219.4800 431.9500 1220.0000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.8500 1219.4800 427.9500 1220.0000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.8500 1219.4800 423.9500 1220.0000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.8500 1219.4800 419.9500 1220.0000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.8500 1219.4800 415.9500 1220.0000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.8500 1219.4800 411.9500 1220.0000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.8500 1219.4800 407.9500 1220.0000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.8500 1219.4800 403.9500 1220.0000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.8500 1219.4800 399.9500 1220.0000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.8500 1219.4800 395.9500 1220.0000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.8500 1219.4800 391.9500 1220.0000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.8500 1219.4800 387.9500 1220.0000 ;
    END
  END out[0]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 643.7500 0.5200 643.8500 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 639.7500 0.5200 639.8500 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 635.7500 0.5200 635.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 631.7500 0.5200 631.8500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 627.7500 0.5200 627.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 623.7500 0.5200 623.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 619.7500 0.5200 619.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 615.7500 0.5200 615.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 611.7500 0.5200 611.8500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 607.7500 0.5200 607.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 603.7500 0.5200 603.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 599.7500 0.5200 599.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 595.7500 0.5200 595.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 591.7500 0.5200 591.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 587.7500 0.5200 587.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 583.7500 0.5200 583.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 579.7500 0.5200 579.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 575.7500 0.5200 575.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 571.7500 0.5200 571.8500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 647.7500 0.5200 647.8500 ;
    END
  END reset
  PIN sum_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.8500 1219.4800 383.9500 1220.0000 ;
    END
  END sum_in[23]
  PIN sum_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.8500 1219.4800 379.9500 1220.0000 ;
    END
  END sum_in[22]
  PIN sum_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.8500 1219.4800 375.9500 1220.0000 ;
    END
  END sum_in[21]
  PIN sum_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.8500 1219.4800 371.9500 1220.0000 ;
    END
  END sum_in[20]
  PIN sum_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.8500 1219.4800 367.9500 1220.0000 ;
    END
  END sum_in[19]
  PIN sum_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.8500 1219.4800 363.9500 1220.0000 ;
    END
  END sum_in[18]
  PIN sum_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.8500 1219.4800 359.9500 1220.0000 ;
    END
  END sum_in[17]
  PIN sum_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.8500 1219.4800 355.9500 1220.0000 ;
    END
  END sum_in[16]
  PIN sum_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.8500 1219.4800 351.9500 1220.0000 ;
    END
  END sum_in[15]
  PIN sum_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.8500 1219.4800 347.9500 1220.0000 ;
    END
  END sum_in[14]
  PIN sum_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.8500 1219.4800 343.9500 1220.0000 ;
    END
  END sum_in[13]
  PIN sum_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.8500 1219.4800 339.9500 1220.0000 ;
    END
  END sum_in[12]
  PIN sum_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.8500 1219.4800 335.9500 1220.0000 ;
    END
  END sum_in[11]
  PIN sum_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.8500 1219.4800 331.9500 1220.0000 ;
    END
  END sum_in[10]
  PIN sum_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.8500 1219.4800 327.9500 1220.0000 ;
    END
  END sum_in[9]
  PIN sum_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.8500 1219.4800 323.9500 1220.0000 ;
    END
  END sum_in[8]
  PIN sum_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.8500 1219.4800 319.9500 1220.0000 ;
    END
  END sum_in[7]
  PIN sum_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.8500 1219.4800 315.9500 1220.0000 ;
    END
  END sum_in[6]
  PIN sum_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.8500 1219.4800 311.9500 1220.0000 ;
    END
  END sum_in[5]
  PIN sum_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.8500 1219.4800 307.9500 1220.0000 ;
    END
  END sum_in[4]
  PIN sum_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.8500 1219.4800 303.9500 1220.0000 ;
    END
  END sum_in[3]
  PIN sum_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.8500 1219.4800 299.9500 1220.0000 ;
    END
  END sum_in[2]
  PIN sum_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.8500 1219.4800 295.9500 1220.0000 ;
    END
  END sum_in[1]
  PIN sum_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.8500 1219.4800 291.9500 1220.0000 ;
    END
  END sum_in[0]
  PIN sfp_sum_fifo_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 651.7500 0.5200 651.8500 ;
    END
  END sfp_sum_fifo_rd
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M5 ;
        RECT 6.0000 303.1800 1214.0000 305.1800 ;
        RECT 6.0000 151.0850 1214.0000 153.0850 ;
        RECT 6.0000 31.0100 1214.0000 33.0100 ;
        RECT 6.0000 23.0050 1214.0000 25.0050 ;
        RECT 6.0000 15.0000 1214.0000 17.0000 ;
        RECT 6.0000 71.0350 1214.0000 73.0350 ;
        RECT 6.0000 63.0300 1214.0000 65.0300 ;
        RECT 6.0000 55.0250 1214.0000 57.0250 ;
        RECT 6.0000 47.0200 1214.0000 49.0200 ;
        RECT 6.0000 39.0150 1214.0000 41.0150 ;
        RECT 6.0000 79.0400 1214.0000 81.0400 ;
        RECT 6.0000 87.0450 1214.0000 89.0450 ;
        RECT 6.0000 95.0500 1214.0000 97.0500 ;
        RECT 6.0000 103.0550 1214.0000 105.0550 ;
        RECT 6.0000 111.0600 1214.0000 113.0600 ;
        RECT 6.0000 119.0650 1214.0000 121.0650 ;
        RECT 6.0000 127.0700 1214.0000 129.0700 ;
        RECT 6.0000 135.0750 1214.0000 137.0750 ;
        RECT 6.0000 143.0800 1214.0000 145.0800 ;
        RECT 6.0000 159.0900 1214.0000 161.0900 ;
        RECT 6.0000 167.0950 1214.0000 169.0950 ;
        RECT 6.0000 175.1000 1214.0000 177.1000 ;
        RECT 6.0000 183.1050 1214.0000 185.1050 ;
        RECT 6.0000 191.1100 1214.0000 193.1100 ;
        RECT 6.0000 199.1150 1214.0000 201.1150 ;
        RECT 6.0000 207.1200 1214.0000 209.1200 ;
        RECT 6.0000 223.1300 1214.0000 225.1300 ;
        RECT 6.0000 215.1250 1214.0000 217.1250 ;
        RECT 6.0000 295.1750 1214.0000 297.1750 ;
        RECT 6.0000 287.1700 1214.0000 289.1700 ;
        RECT 6.0000 279.1650 1214.0000 281.1650 ;
        RECT 6.0000 271.1600 1214.0000 273.1600 ;
        RECT 6.0000 263.1550 1214.0000 265.1550 ;
        RECT 6.0000 255.1500 1214.0000 257.1500 ;
        RECT 6.0000 247.1450 1214.0000 249.1450 ;
        RECT 6.0000 239.1400 1214.0000 241.1400 ;
        RECT 6.0000 231.1350 1214.0000 233.1350 ;
        RECT 6.0000 311.1850 1214.0000 313.1850 ;
        RECT 6.0000 335.2000 1214.0000 337.2000 ;
        RECT 6.0000 327.1950 1214.0000 329.1950 ;
        RECT 6.0000 319.1900 1214.0000 321.1900 ;
        RECT 6.0000 343.2050 1214.0000 345.2050 ;
        RECT 6.0000 351.2100 1214.0000 353.2100 ;
        RECT 6.0000 359.2150 1214.0000 361.2150 ;
        RECT 6.0000 367.2200 1214.0000 369.2200 ;
        RECT 6.0000 375.2250 1214.0000 377.2250 ;
        RECT 6.0000 399.2400 1214.0000 401.2400 ;
        RECT 6.0000 391.2350 1214.0000 393.2350 ;
        RECT 6.0000 383.2300 1214.0000 385.2300 ;
        RECT 6.0000 415.2500 1214.0000 417.2500 ;
        RECT 6.0000 407.2450 1214.0000 409.2450 ;
        RECT 6.0000 431.2600 1214.0000 433.2600 ;
        RECT 6.0000 423.2550 1214.0000 425.2550 ;
        RECT 6.0000 455.2750 1214.0000 457.2750 ;
        RECT 6.0000 447.2700 1214.0000 449.2700 ;
        RECT 6.0000 439.2650 1214.0000 441.2650 ;
        RECT 6.0000 495.3000 1214.0000 497.3000 ;
        RECT 6.0000 471.2850 1214.0000 473.2850 ;
        RECT 6.0000 463.2800 1214.0000 465.2800 ;
        RECT 6.0000 479.2900 1214.0000 481.2900 ;
        RECT 6.0000 487.2950 1214.0000 489.2950 ;
        RECT 6.0000 527.3200 1214.0000 529.3200 ;
        RECT 6.0000 519.3150 1214.0000 521.3150 ;
        RECT 6.0000 511.3100 1214.0000 513.3100 ;
        RECT 6.0000 503.3050 1214.0000 505.3050 ;
        RECT 6.0000 535.3250 1214.0000 537.3250 ;
        RECT 6.0000 543.3300 1214.0000 545.3300 ;
        RECT 6.0000 551.3350 1214.0000 553.3350 ;
        RECT 6.0000 559.3400 1214.0000 561.3400 ;
        RECT 6.0000 567.3450 1214.0000 569.3450 ;
        RECT 6.0000 575.3500 1214.0000 577.3500 ;
        RECT 6.0000 583.3550 1214.0000 585.3550 ;
        RECT 6.0000 591.3600 1214.0000 593.3600 ;
        RECT 6.0000 599.3650 1214.0000 601.3650 ;
        RECT 6.0000 607.3700 1214.0000 609.3700 ;
        RECT 6.0000 615.3750 1214.0000 617.3750 ;
        RECT 6.0000 623.3800 1214.0000 625.3800 ;
        RECT 6.0000 631.3850 1214.0000 633.3850 ;
        RECT 6.0000 639.3900 1214.0000 641.3900 ;
        RECT 6.0000 647.3950 1214.0000 649.3950 ;
        RECT 6.0000 655.4000 1214.0000 657.4000 ;
        RECT 6.0000 663.4050 1214.0000 665.4050 ;
        RECT 6.0000 671.4100 1214.0000 673.4100 ;
        RECT 6.0000 679.4150 1214.0000 681.4150 ;
        RECT 6.0000 759.4650 1214.0000 761.4650 ;
        RECT 6.0000 751.4600 1214.0000 753.4600 ;
        RECT 6.0000 743.4550 1214.0000 745.4550 ;
        RECT 6.0000 735.4500 1214.0000 737.4500 ;
        RECT 6.0000 727.4450 1214.0000 729.4450 ;
        RECT 6.0000 719.4400 1214.0000 721.4400 ;
        RECT 6.0000 711.4350 1214.0000 713.4350 ;
        RECT 6.0000 703.4300 1214.0000 705.4300 ;
        RECT 6.0000 695.4250 1214.0000 697.4250 ;
        RECT 6.0000 687.4200 1214.0000 689.4200 ;
        RECT 6.0000 767.4700 1214.0000 769.4700 ;
        RECT 6.0000 775.4750 1214.0000 777.4750 ;
        RECT 6.0000 783.4800 1214.0000 785.4800 ;
        RECT 6.0000 791.4850 1214.0000 793.4850 ;
        RECT 6.0000 799.4900 1214.0000 801.4900 ;
        RECT 6.0000 807.4950 1214.0000 809.4950 ;
        RECT 6.0000 815.5000 1214.0000 817.5000 ;
        RECT 6.0000 831.5100 1214.0000 833.5100 ;
        RECT 6.0000 823.5050 1214.0000 825.5050 ;
        RECT 6.0000 911.5600 1214.0000 913.5600 ;
        RECT 6.0000 903.5550 1214.0000 905.5550 ;
        RECT 6.0000 895.5500 1214.0000 897.5500 ;
        RECT 6.0000 887.5450 1214.0000 889.5450 ;
        RECT 6.0000 879.5400 1214.0000 881.5400 ;
        RECT 6.0000 871.5350 1214.0000 873.5350 ;
        RECT 6.0000 863.5300 1214.0000 865.5300 ;
        RECT 6.0000 855.5250 1214.0000 857.5250 ;
        RECT 6.0000 847.5200 1214.0000 849.5200 ;
        RECT 6.0000 839.5150 1214.0000 841.5150 ;
        RECT 6.0000 919.5650 1214.0000 921.5650 ;
        RECT 6.0000 927.5700 1214.0000 929.5700 ;
        RECT 6.0000 935.5750 1214.0000 937.5750 ;
        RECT 6.0000 943.5800 1214.0000 945.5800 ;
        RECT 6.0000 951.5850 1214.0000 953.5850 ;
        RECT 6.0000 959.5900 1214.0000 961.5900 ;
        RECT 6.0000 967.5950 1214.0000 969.5950 ;
        RECT 6.0000 983.6050 1214.0000 985.6050 ;
        RECT 6.0000 975.6000 1214.0000 977.6000 ;
        RECT 6.0000 1063.6550 1214.0000 1065.6550 ;
        RECT 6.0000 1055.6500 1214.0000 1057.6500 ;
        RECT 6.0000 1047.6450 1214.0000 1049.6450 ;
        RECT 6.0000 1039.6400 1214.0000 1041.6400 ;
        RECT 6.0000 1031.6350 1214.0000 1033.6350 ;
        RECT 6.0000 1023.6300 1214.0000 1025.6300 ;
        RECT 6.0000 1015.6250 1214.0000 1017.6250 ;
        RECT 6.0000 1007.6200 1214.0000 1009.6200 ;
        RECT 6.0000 999.6150 1214.0000 1001.6150 ;
        RECT 6.0000 991.6100 1214.0000 993.6100 ;
        RECT 6.0000 1143.7050 1214.0000 1145.7050 ;
        RECT 6.0000 1071.6600 1214.0000 1073.6600 ;
        RECT 6.0000 1079.6650 1214.0000 1081.6650 ;
        RECT 6.0000 1087.6700 1214.0000 1089.6700 ;
        RECT 6.0000 1095.6750 1214.0000 1097.6750 ;
        RECT 6.0000 1103.6800 1214.0000 1105.6800 ;
        RECT 6.0000 1111.6850 1214.0000 1113.6850 ;
        RECT 6.0000 1119.6900 1214.0000 1121.6900 ;
        RECT 6.0000 1127.6950 1214.0000 1129.6950 ;
        RECT 6.0000 1135.7000 1214.0000 1137.7000 ;
        RECT 6.0000 1175.7250 1214.0000 1177.7250 ;
        RECT 6.0000 1167.7200 1214.0000 1169.7200 ;
        RECT 6.0000 1159.7150 1214.0000 1161.7150 ;
        RECT 6.0000 1151.7100 1214.0000 1153.7100 ;
        RECT 6.0000 1207.7450 1214.0000 1209.7450 ;
        RECT 6.0000 1199.7400 1214.0000 1201.7400 ;
        RECT 6.0000 1191.7350 1214.0000 1193.7350 ;
        RECT 6.0000 1183.7300 1214.0000 1185.7300 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M5 ;
        RECT 2.0000 10.0000 1218.0000 12.0000 ;
        RECT 2.0000 18.0050 1218.0000 20.0050 ;
        RECT 2.0000 26.0100 1218.0000 28.0100 ;
        RECT 2.0000 34.0150 1218.0000 36.0150 ;
        RECT 2.0000 42.0200 1218.0000 44.0200 ;
        RECT 2.0000 50.0250 1218.0000 52.0250 ;
        RECT 2.0000 58.0300 1218.0000 60.0300 ;
        RECT 2.0000 74.0400 1218.0000 76.0400 ;
        RECT 2.0000 66.0350 1218.0000 68.0350 ;
        RECT 2.0000 82.0450 1218.0000 84.0450 ;
        RECT 2.0000 90.0500 1218.0000 92.0500 ;
        RECT 2.0000 98.0550 1218.0000 100.0550 ;
        RECT 2.0000 106.0600 1218.0000 108.0600 ;
        RECT 2.0000 114.0650 1218.0000 116.0650 ;
        RECT 2.0000 122.0700 1218.0000 124.0700 ;
        RECT 2.0000 130.0750 1218.0000 132.0750 ;
        RECT 2.0000 138.0800 1218.0000 140.0800 ;
        RECT 2.0000 146.0850 1218.0000 148.0850 ;
        RECT 2.0000 154.0900 1218.0000 156.0900 ;
        RECT 2.0000 162.0950 1218.0000 164.0950 ;
        RECT 2.0000 170.1000 1218.0000 172.1000 ;
        RECT 2.0000 178.1050 1218.0000 180.1050 ;
        RECT 2.0000 186.1100 1218.0000 188.1100 ;
        RECT 2.0000 194.1150 1218.0000 196.1150 ;
        RECT 2.0000 202.1200 1218.0000 204.1200 ;
        RECT 2.0000 210.1250 1218.0000 212.1250 ;
        RECT 2.0000 218.1300 1218.0000 220.1300 ;
        RECT 2.0000 226.1350 1218.0000 228.1350 ;
        RECT 2.0000 234.1400 1218.0000 236.1400 ;
        RECT 2.0000 242.1450 1218.0000 244.1450 ;
        RECT 2.0000 250.1500 1218.0000 252.1500 ;
        RECT 2.0000 258.1550 1218.0000 260.1550 ;
        RECT 2.0000 266.1600 1218.0000 268.1600 ;
        RECT 2.0000 274.1650 1218.0000 276.1650 ;
        RECT 2.0000 282.1700 1218.0000 284.1700 ;
        RECT 2.0000 290.1750 1218.0000 292.1750 ;
        RECT 2.0000 298.1800 1218.0000 300.1800 ;
        RECT 2.0000 306.1850 1218.0000 308.1850 ;
        RECT 2.0000 314.1900 1218.0000 316.1900 ;
        RECT 2.0000 322.1950 1218.0000 324.1950 ;
        RECT 2.0000 330.2000 1218.0000 332.2000 ;
        RECT 2.0000 338.2050 1218.0000 340.2050 ;
        RECT 2.0000 354.2150 1218.0000 356.2150 ;
        RECT 2.0000 346.2100 1218.0000 348.2100 ;
        RECT 2.0000 362.2200 1218.0000 364.2200 ;
        RECT 2.0000 378.2300 1218.0000 380.2300 ;
        RECT 2.0000 370.2250 1218.0000 372.2250 ;
        RECT 2.0000 418.2550 1218.0000 420.2550 ;
        RECT 2.0000 394.2400 1218.0000 396.2400 ;
        RECT 2.0000 386.2350 1218.0000 388.2350 ;
        RECT 2.0000 410.2500 1218.0000 412.2500 ;
        RECT 2.0000 402.2450 1218.0000 404.2450 ;
        RECT 2.0000 434.2650 1218.0000 436.2650 ;
        RECT 2.0000 426.2600 1218.0000 428.2600 ;
        RECT 2.0000 450.2750 1218.0000 452.2750 ;
        RECT 2.0000 442.2700 1218.0000 444.2700 ;
        RECT 2.0000 474.2900 1218.0000 476.2900 ;
        RECT 2.0000 466.2850 1218.0000 468.2850 ;
        RECT 2.0000 458.2800 1218.0000 460.2800 ;
        RECT 2.0000 490.3000 1218.0000 492.3000 ;
        RECT 2.0000 482.2950 1218.0000 484.2950 ;
        RECT 2.0000 498.3050 1218.0000 500.3050 ;
        RECT 2.0000 506.3100 1218.0000 508.3100 ;
        RECT 2.0000 514.3150 1218.0000 516.3150 ;
        RECT 2.0000 522.3200 1218.0000 524.3200 ;
        RECT 2.0000 530.3250 1218.0000 532.3250 ;
        RECT 2.0000 602.3700 1218.0000 604.3700 ;
        RECT 2.0000 594.3650 1218.0000 596.3650 ;
        RECT 2.0000 586.3600 1218.0000 588.3600 ;
        RECT 2.0000 578.3550 1218.0000 580.3550 ;
        RECT 2.0000 570.3500 1218.0000 572.3500 ;
        RECT 2.0000 562.3450 1218.0000 564.3450 ;
        RECT 2.0000 554.3400 1218.0000 556.3400 ;
        RECT 2.0000 546.3350 1218.0000 548.3350 ;
        RECT 2.0000 538.3300 1218.0000 540.3300 ;
        RECT 2.0000 914.5650 1218.0000 916.5650 ;
        RECT 2.0000 762.4700 1218.0000 764.4700 ;
        RECT 2.0000 674.4150 1218.0000 676.4150 ;
        RECT 2.0000 682.4200 1218.0000 684.4200 ;
        RECT 2.0000 666.4100 1218.0000 668.4100 ;
        RECT 2.0000 658.4050 1218.0000 660.4050 ;
        RECT 2.0000 650.4000 1218.0000 652.4000 ;
        RECT 2.0000 642.3950 1218.0000 644.3950 ;
        RECT 2.0000 634.3900 1218.0000 636.3900 ;
        RECT 2.0000 626.3850 1218.0000 628.3850 ;
        RECT 2.0000 618.3800 1218.0000 620.3800 ;
        RECT 2.0000 610.3750 1218.0000 612.3750 ;
        RECT 2.0000 690.4250 1218.0000 692.4250 ;
        RECT 2.0000 698.4300 1218.0000 700.4300 ;
        RECT 2.0000 706.4350 1218.0000 708.4350 ;
        RECT 2.0000 714.4400 1218.0000 716.4400 ;
        RECT 2.0000 722.4450 1218.0000 724.4450 ;
        RECT 2.0000 730.4500 1218.0000 732.4500 ;
        RECT 2.0000 738.4550 1218.0000 740.4550 ;
        RECT 2.0000 746.4600 1218.0000 748.4600 ;
        RECT 2.0000 754.4650 1218.0000 756.4650 ;
        RECT 2.0000 770.4750 1218.0000 772.4750 ;
        RECT 2.0000 778.4800 1218.0000 780.4800 ;
        RECT 2.0000 786.4850 1218.0000 788.4850 ;
        RECT 2.0000 794.4900 1218.0000 796.4900 ;
        RECT 2.0000 802.4950 1218.0000 804.4950 ;
        RECT 2.0000 810.5000 1218.0000 812.5000 ;
        RECT 2.0000 818.5050 1218.0000 820.5050 ;
        RECT 2.0000 826.5100 1218.0000 828.5100 ;
        RECT 2.0000 834.5150 1218.0000 836.5150 ;
        RECT 2.0000 842.5200 1218.0000 844.5200 ;
        RECT 2.0000 850.5250 1218.0000 852.5250 ;
        RECT 2.0000 858.5300 1218.0000 860.5300 ;
        RECT 2.0000 866.5350 1218.0000 868.5350 ;
        RECT 2.0000 874.5400 1218.0000 876.5400 ;
        RECT 2.0000 882.5450 1218.0000 884.5450 ;
        RECT 2.0000 890.5500 1218.0000 892.5500 ;
        RECT 2.0000 898.5550 1218.0000 900.5550 ;
        RECT 2.0000 906.5600 1218.0000 908.5600 ;
        RECT 2.0000 1066.6600 1218.0000 1068.6600 ;
        RECT 2.0000 962.5950 1218.0000 964.5950 ;
        RECT 2.0000 986.6100 1218.0000 988.6100 ;
        RECT 2.0000 978.6050 1218.0000 980.6050 ;
        RECT 2.0000 970.6000 1218.0000 972.6000 ;
        RECT 2.0000 954.5900 1218.0000 956.5900 ;
        RECT 2.0000 946.5850 1218.0000 948.5850 ;
        RECT 2.0000 938.5800 1218.0000 940.5800 ;
        RECT 2.0000 930.5750 1218.0000 932.5750 ;
        RECT 2.0000 922.5700 1218.0000 924.5700 ;
        RECT 2.0000 1058.6550 1218.0000 1060.6550 ;
        RECT 2.0000 1050.6500 1218.0000 1052.6500 ;
        RECT 2.0000 1042.6450 1218.0000 1044.6450 ;
        RECT 2.0000 1034.6400 1218.0000 1036.6400 ;
        RECT 2.0000 1026.6350 1218.0000 1028.6350 ;
        RECT 2.0000 1018.6300 1218.0000 1020.6300 ;
        RECT 2.0000 1010.6250 1218.0000 1012.6250 ;
        RECT 2.0000 1002.6200 1218.0000 1004.6200 ;
        RECT 2.0000 994.6150 1218.0000 996.6150 ;
        RECT 2.0000 1138.7050 1218.0000 1140.7050 ;
        RECT 2.0000 1130.7000 1218.0000 1132.7000 ;
        RECT 2.0000 1122.6950 1218.0000 1124.6950 ;
        RECT 2.0000 1114.6900 1218.0000 1116.6900 ;
        RECT 2.0000 1106.6850 1218.0000 1108.6850 ;
        RECT 2.0000 1098.6800 1218.0000 1100.6800 ;
        RECT 2.0000 1090.6750 1218.0000 1092.6750 ;
        RECT 2.0000 1082.6700 1218.0000 1084.6700 ;
        RECT 2.0000 1074.6650 1218.0000 1076.6650 ;
        RECT 2.0000 1146.7100 1218.0000 1148.7100 ;
        RECT 2.0000 1154.7150 1218.0000 1156.7150 ;
        RECT 2.0000 1162.7200 1218.0000 1164.7200 ;
        RECT 2.0000 1170.7250 1218.0000 1172.7250 ;
        RECT 2.0000 1178.7300 1218.0000 1180.7300 ;
        RECT 2.0000 1186.7350 1218.0000 1188.7350 ;
        RECT 2.0000 1194.7400 1218.0000 1196.7400 ;
        RECT 2.0000 1202.7450 1218.0000 1204.7450 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1220.0000 1220.0000 ;
    LAYER M2 ;
      RECT 1024.0500 1219.3800 1220.0000 1220.0000 ;
      RECT 1020.0500 1219.3800 1023.7500 1220.0000 ;
      RECT 1016.0500 1219.3800 1019.7500 1220.0000 ;
      RECT 1012.0500 1219.3800 1015.7500 1220.0000 ;
      RECT 1008.0500 1219.3800 1011.7500 1220.0000 ;
      RECT 1004.0500 1219.3800 1007.7500 1220.0000 ;
      RECT 1000.0500 1219.3800 1003.7500 1220.0000 ;
      RECT 996.0500 1219.3800 999.7500 1220.0000 ;
      RECT 992.0500 1219.3800 995.7500 1220.0000 ;
      RECT 988.0500 1219.3800 991.7500 1220.0000 ;
      RECT 984.0500 1219.3800 987.7500 1220.0000 ;
      RECT 980.0500 1219.3800 983.7500 1220.0000 ;
      RECT 976.0500 1219.3800 979.7500 1220.0000 ;
      RECT 972.0500 1219.3800 975.7500 1220.0000 ;
      RECT 968.0500 1219.3800 971.7500 1220.0000 ;
      RECT 964.0500 1219.3800 967.7500 1220.0000 ;
      RECT 960.0500 1219.3800 963.7500 1220.0000 ;
      RECT 956.0500 1219.3800 959.7500 1220.0000 ;
      RECT 952.0500 1219.3800 955.7500 1220.0000 ;
      RECT 948.0500 1219.3800 951.7500 1220.0000 ;
      RECT 944.0500 1219.3800 947.7500 1220.0000 ;
      RECT 940.0500 1219.3800 943.7500 1220.0000 ;
      RECT 936.0500 1219.3800 939.7500 1220.0000 ;
      RECT 932.0500 1219.3800 935.7500 1220.0000 ;
      RECT 928.0500 1219.3800 931.7500 1220.0000 ;
      RECT 924.0500 1219.3800 927.7500 1220.0000 ;
      RECT 920.0500 1219.3800 923.7500 1220.0000 ;
      RECT 916.0500 1219.3800 919.7500 1220.0000 ;
      RECT 912.0500 1219.3800 915.7500 1220.0000 ;
      RECT 908.0500 1219.3800 911.7500 1220.0000 ;
      RECT 904.0500 1219.3800 907.7500 1220.0000 ;
      RECT 900.0500 1219.3800 903.7500 1220.0000 ;
      RECT 896.0500 1219.3800 899.7500 1220.0000 ;
      RECT 892.0500 1219.3800 895.7500 1220.0000 ;
      RECT 888.0500 1219.3800 891.7500 1220.0000 ;
      RECT 884.0500 1219.3800 887.7500 1220.0000 ;
      RECT 880.0500 1219.3800 883.7500 1220.0000 ;
      RECT 876.0500 1219.3800 879.7500 1220.0000 ;
      RECT 872.0500 1219.3800 875.7500 1220.0000 ;
      RECT 868.0500 1219.3800 871.7500 1220.0000 ;
      RECT 864.0500 1219.3800 867.7500 1220.0000 ;
      RECT 860.0500 1219.3800 863.7500 1220.0000 ;
      RECT 856.0500 1219.3800 859.7500 1220.0000 ;
      RECT 852.0500 1219.3800 855.7500 1220.0000 ;
      RECT 848.0500 1219.3800 851.7500 1220.0000 ;
      RECT 844.0500 1219.3800 847.7500 1220.0000 ;
      RECT 840.0500 1219.3800 843.7500 1220.0000 ;
      RECT 836.0500 1219.3800 839.7500 1220.0000 ;
      RECT 832.0500 1219.3800 835.7500 1220.0000 ;
      RECT 828.0500 1219.3800 831.7500 1220.0000 ;
      RECT 824.0500 1219.3800 827.7500 1220.0000 ;
      RECT 820.0500 1219.3800 823.7500 1220.0000 ;
      RECT 816.0500 1219.3800 819.7500 1220.0000 ;
      RECT 812.0500 1219.3800 815.7500 1220.0000 ;
      RECT 808.0500 1219.3800 811.7500 1220.0000 ;
      RECT 804.0500 1219.3800 807.7500 1220.0000 ;
      RECT 800.0500 1219.3800 803.7500 1220.0000 ;
      RECT 796.0500 1219.3800 799.7500 1220.0000 ;
      RECT 792.0500 1219.3800 795.7500 1220.0000 ;
      RECT 788.0500 1219.3800 791.7500 1220.0000 ;
      RECT 784.0500 1219.3800 787.7500 1220.0000 ;
      RECT 780.0500 1219.3800 783.7500 1220.0000 ;
      RECT 776.0500 1219.3800 779.7500 1220.0000 ;
      RECT 772.0500 1219.3800 775.7500 1220.0000 ;
      RECT 768.0500 1219.3800 771.7500 1220.0000 ;
      RECT 764.0500 1219.3800 767.7500 1220.0000 ;
      RECT 760.0500 1219.3800 763.7500 1220.0000 ;
      RECT 756.0500 1219.3800 759.7500 1220.0000 ;
      RECT 752.0500 1219.3800 755.7500 1220.0000 ;
      RECT 748.0500 1219.3800 751.7500 1220.0000 ;
      RECT 744.0500 1219.3800 747.7500 1220.0000 ;
      RECT 740.0500 1219.3800 743.7500 1220.0000 ;
      RECT 736.0500 1219.3800 739.7500 1220.0000 ;
      RECT 732.0500 1219.3800 735.7500 1220.0000 ;
      RECT 728.0500 1219.3800 731.7500 1220.0000 ;
      RECT 724.0500 1219.3800 727.7500 1220.0000 ;
      RECT 720.0500 1219.3800 723.7500 1220.0000 ;
      RECT 716.0500 1219.3800 719.7500 1220.0000 ;
      RECT 712.0500 1219.3800 715.7500 1220.0000 ;
      RECT 708.0500 1219.3800 711.7500 1220.0000 ;
      RECT 704.0500 1219.3800 707.7500 1220.0000 ;
      RECT 700.0500 1219.3800 703.7500 1220.0000 ;
      RECT 696.0500 1219.3800 699.7500 1220.0000 ;
      RECT 692.0500 1219.3800 695.7500 1220.0000 ;
      RECT 688.0500 1219.3800 691.7500 1220.0000 ;
      RECT 684.0500 1219.3800 687.7500 1220.0000 ;
      RECT 680.0500 1219.3800 683.7500 1220.0000 ;
      RECT 676.0500 1219.3800 679.7500 1220.0000 ;
      RECT 672.0500 1219.3800 675.7500 1220.0000 ;
      RECT 668.0500 1219.3800 671.7500 1220.0000 ;
      RECT 664.0500 1219.3800 667.7500 1220.0000 ;
      RECT 660.0500 1219.3800 663.7500 1220.0000 ;
      RECT 656.0500 1219.3800 659.7500 1220.0000 ;
      RECT 652.0500 1219.3800 655.7500 1220.0000 ;
      RECT 648.0500 1219.3800 651.7500 1220.0000 ;
      RECT 644.0500 1219.3800 647.7500 1220.0000 ;
      RECT 640.0500 1219.3800 643.7500 1220.0000 ;
      RECT 636.0500 1219.3800 639.7500 1220.0000 ;
      RECT 632.0500 1219.3800 635.7500 1220.0000 ;
      RECT 628.0500 1219.3800 631.7500 1220.0000 ;
      RECT 624.0500 1219.3800 627.7500 1220.0000 ;
      RECT 620.0500 1219.3800 623.7500 1220.0000 ;
      RECT 616.0500 1219.3800 619.7500 1220.0000 ;
      RECT 612.0500 1219.3800 615.7500 1220.0000 ;
      RECT 608.0500 1219.3800 611.7500 1220.0000 ;
      RECT 604.0500 1219.3800 607.7500 1220.0000 ;
      RECT 600.0500 1219.3800 603.7500 1220.0000 ;
      RECT 596.0500 1219.3800 599.7500 1220.0000 ;
      RECT 592.0500 1219.3800 595.7500 1220.0000 ;
      RECT 588.0500 1219.3800 591.7500 1220.0000 ;
      RECT 584.0500 1219.3800 587.7500 1220.0000 ;
      RECT 580.0500 1219.3800 583.7500 1220.0000 ;
      RECT 576.0500 1219.3800 579.7500 1220.0000 ;
      RECT 572.0500 1219.3800 575.7500 1220.0000 ;
      RECT 568.0500 1219.3800 571.7500 1220.0000 ;
      RECT 564.0500 1219.3800 567.7500 1220.0000 ;
      RECT 560.0500 1219.3800 563.7500 1220.0000 ;
      RECT 556.0500 1219.3800 559.7500 1220.0000 ;
      RECT 552.0500 1219.3800 555.7500 1220.0000 ;
      RECT 548.0500 1219.3800 551.7500 1220.0000 ;
      RECT 544.0500 1219.3800 547.7500 1220.0000 ;
      RECT 540.0500 1219.3800 543.7500 1220.0000 ;
      RECT 536.0500 1219.3800 539.7500 1220.0000 ;
      RECT 532.0500 1219.3800 535.7500 1220.0000 ;
      RECT 528.0500 1219.3800 531.7500 1220.0000 ;
      RECT 524.0500 1219.3800 527.7500 1220.0000 ;
      RECT 520.0500 1219.3800 523.7500 1220.0000 ;
      RECT 516.0500 1219.3800 519.7500 1220.0000 ;
      RECT 512.0500 1219.3800 515.7500 1220.0000 ;
      RECT 508.0500 1219.3800 511.7500 1220.0000 ;
      RECT 504.0500 1219.3800 507.7500 1220.0000 ;
      RECT 500.0500 1219.3800 503.7500 1220.0000 ;
      RECT 496.0500 1219.3800 499.7500 1220.0000 ;
      RECT 492.0500 1219.3800 495.7500 1220.0000 ;
      RECT 488.0500 1219.3800 491.7500 1220.0000 ;
      RECT 484.0500 1219.3800 487.7500 1220.0000 ;
      RECT 480.0500 1219.3800 483.7500 1220.0000 ;
      RECT 476.0500 1219.3800 479.7500 1220.0000 ;
      RECT 472.0500 1219.3800 475.7500 1220.0000 ;
      RECT 468.0500 1219.3800 471.7500 1220.0000 ;
      RECT 464.0500 1219.3800 467.7500 1220.0000 ;
      RECT 460.0500 1219.3800 463.7500 1220.0000 ;
      RECT 456.0500 1219.3800 459.7500 1220.0000 ;
      RECT 452.0500 1219.3800 455.7500 1220.0000 ;
      RECT 448.0500 1219.3800 451.7500 1220.0000 ;
      RECT 444.0500 1219.3800 447.7500 1220.0000 ;
      RECT 440.0500 1219.3800 443.7500 1220.0000 ;
      RECT 436.0500 1219.3800 439.7500 1220.0000 ;
      RECT 432.0500 1219.3800 435.7500 1220.0000 ;
      RECT 428.0500 1219.3800 431.7500 1220.0000 ;
      RECT 424.0500 1219.3800 427.7500 1220.0000 ;
      RECT 420.0500 1219.3800 423.7500 1220.0000 ;
      RECT 416.0500 1219.3800 419.7500 1220.0000 ;
      RECT 412.0500 1219.3800 415.7500 1220.0000 ;
      RECT 408.0500 1219.3800 411.7500 1220.0000 ;
      RECT 404.0500 1219.3800 407.7500 1220.0000 ;
      RECT 400.0500 1219.3800 403.7500 1220.0000 ;
      RECT 396.0500 1219.3800 399.7500 1220.0000 ;
      RECT 392.0500 1219.3800 395.7500 1220.0000 ;
      RECT 388.0500 1219.3800 391.7500 1220.0000 ;
      RECT 384.0500 1219.3800 387.7500 1220.0000 ;
      RECT 380.0500 1219.3800 383.7500 1220.0000 ;
      RECT 376.0500 1219.3800 379.7500 1220.0000 ;
      RECT 372.0500 1219.3800 375.7500 1220.0000 ;
      RECT 368.0500 1219.3800 371.7500 1220.0000 ;
      RECT 364.0500 1219.3800 367.7500 1220.0000 ;
      RECT 360.0500 1219.3800 363.7500 1220.0000 ;
      RECT 356.0500 1219.3800 359.7500 1220.0000 ;
      RECT 352.0500 1219.3800 355.7500 1220.0000 ;
      RECT 348.0500 1219.3800 351.7500 1220.0000 ;
      RECT 344.0500 1219.3800 347.7500 1220.0000 ;
      RECT 340.0500 1219.3800 343.7500 1220.0000 ;
      RECT 336.0500 1219.3800 339.7500 1220.0000 ;
      RECT 332.0500 1219.3800 335.7500 1220.0000 ;
      RECT 328.0500 1219.3800 331.7500 1220.0000 ;
      RECT 324.0500 1219.3800 327.7500 1220.0000 ;
      RECT 320.0500 1219.3800 323.7500 1220.0000 ;
      RECT 316.0500 1219.3800 319.7500 1220.0000 ;
      RECT 312.0500 1219.3800 315.7500 1220.0000 ;
      RECT 308.0500 1219.3800 311.7500 1220.0000 ;
      RECT 304.0500 1219.3800 307.7500 1220.0000 ;
      RECT 300.0500 1219.3800 303.7500 1220.0000 ;
      RECT 296.0500 1219.3800 299.7500 1220.0000 ;
      RECT 292.0500 1219.3800 295.7500 1220.0000 ;
      RECT 288.0500 1219.3800 291.7500 1220.0000 ;
      RECT 284.0500 1219.3800 287.7500 1220.0000 ;
      RECT 280.0500 1219.3800 283.7500 1220.0000 ;
      RECT 276.0500 1219.3800 279.7500 1220.0000 ;
      RECT 272.0500 1219.3800 275.7500 1220.0000 ;
      RECT 268.0500 1219.3800 271.7500 1220.0000 ;
      RECT 264.0500 1219.3800 267.7500 1220.0000 ;
      RECT 260.0500 1219.3800 263.7500 1220.0000 ;
      RECT 256.0500 1219.3800 259.7500 1220.0000 ;
      RECT 252.0500 1219.3800 255.7500 1220.0000 ;
      RECT 248.0500 1219.3800 251.7500 1220.0000 ;
      RECT 244.0500 1219.3800 247.7500 1220.0000 ;
      RECT 240.0500 1219.3800 243.7500 1220.0000 ;
      RECT 236.0500 1219.3800 239.7500 1220.0000 ;
      RECT 232.0500 1219.3800 235.7500 1220.0000 ;
      RECT 228.0500 1219.3800 231.7500 1220.0000 ;
      RECT 224.0500 1219.3800 227.7500 1220.0000 ;
      RECT 220.0500 1219.3800 223.7500 1220.0000 ;
      RECT 216.0500 1219.3800 219.7500 1220.0000 ;
      RECT 212.0500 1219.3800 215.7500 1220.0000 ;
      RECT 208.0500 1219.3800 211.7500 1220.0000 ;
      RECT 204.0500 1219.3800 207.7500 1220.0000 ;
      RECT 200.0500 1219.3800 203.7500 1220.0000 ;
      RECT 196.0500 1219.3800 199.7500 1220.0000 ;
      RECT 0.0000 1219.3800 195.7500 1220.0000 ;
      RECT 0.0000 0.6200 1220.0000 1219.3800 ;
      RECT 736.0500 0.0000 1220.0000 0.6200 ;
      RECT 732.0500 0.0000 735.7500 0.6200 ;
      RECT 728.0500 0.0000 731.7500 0.6200 ;
      RECT 724.0500 0.0000 727.7500 0.6200 ;
      RECT 720.0500 0.0000 723.7500 0.6200 ;
      RECT 716.0500 0.0000 719.7500 0.6200 ;
      RECT 712.0500 0.0000 715.7500 0.6200 ;
      RECT 708.0500 0.0000 711.7500 0.6200 ;
      RECT 704.0500 0.0000 707.7500 0.6200 ;
      RECT 700.0500 0.0000 703.7500 0.6200 ;
      RECT 696.0500 0.0000 699.7500 0.6200 ;
      RECT 692.0500 0.0000 695.7500 0.6200 ;
      RECT 688.0500 0.0000 691.7500 0.6200 ;
      RECT 684.0500 0.0000 687.7500 0.6200 ;
      RECT 680.0500 0.0000 683.7500 0.6200 ;
      RECT 676.0500 0.0000 679.7500 0.6200 ;
      RECT 672.0500 0.0000 675.7500 0.6200 ;
      RECT 668.0500 0.0000 671.7500 0.6200 ;
      RECT 664.0500 0.0000 667.7500 0.6200 ;
      RECT 660.0500 0.0000 663.7500 0.6200 ;
      RECT 656.0500 0.0000 659.7500 0.6200 ;
      RECT 652.0500 0.0000 655.7500 0.6200 ;
      RECT 648.0500 0.0000 651.7500 0.6200 ;
      RECT 644.0500 0.0000 647.7500 0.6200 ;
      RECT 640.0500 0.0000 643.7500 0.6200 ;
      RECT 636.0500 0.0000 639.7500 0.6200 ;
      RECT 632.0500 0.0000 635.7500 0.6200 ;
      RECT 628.0500 0.0000 631.7500 0.6200 ;
      RECT 624.0500 0.0000 627.7500 0.6200 ;
      RECT 620.0500 0.0000 623.7500 0.6200 ;
      RECT 616.0500 0.0000 619.7500 0.6200 ;
      RECT 612.0500 0.0000 615.7500 0.6200 ;
      RECT 608.0500 0.0000 611.7500 0.6200 ;
      RECT 604.0500 0.0000 607.7500 0.6200 ;
      RECT 600.0500 0.0000 603.7500 0.6200 ;
      RECT 596.0500 0.0000 599.7500 0.6200 ;
      RECT 592.0500 0.0000 595.7500 0.6200 ;
      RECT 588.0500 0.0000 591.7500 0.6200 ;
      RECT 584.0500 0.0000 587.7500 0.6200 ;
      RECT 580.0500 0.0000 583.7500 0.6200 ;
      RECT 576.0500 0.0000 579.7500 0.6200 ;
      RECT 572.0500 0.0000 575.7500 0.6200 ;
      RECT 568.0500 0.0000 571.7500 0.6200 ;
      RECT 564.0500 0.0000 567.7500 0.6200 ;
      RECT 560.0500 0.0000 563.7500 0.6200 ;
      RECT 556.0500 0.0000 559.7500 0.6200 ;
      RECT 552.0500 0.0000 555.7500 0.6200 ;
      RECT 548.0500 0.0000 551.7500 0.6200 ;
      RECT 544.0500 0.0000 547.7500 0.6200 ;
      RECT 540.0500 0.0000 543.7500 0.6200 ;
      RECT 536.0500 0.0000 539.7500 0.6200 ;
      RECT 532.0500 0.0000 535.7500 0.6200 ;
      RECT 528.0500 0.0000 531.7500 0.6200 ;
      RECT 524.0500 0.0000 527.7500 0.6200 ;
      RECT 520.0500 0.0000 523.7500 0.6200 ;
      RECT 516.0500 0.0000 519.7500 0.6200 ;
      RECT 512.0500 0.0000 515.7500 0.6200 ;
      RECT 508.0500 0.0000 511.7500 0.6200 ;
      RECT 504.0500 0.0000 507.7500 0.6200 ;
      RECT 500.0500 0.0000 503.7500 0.6200 ;
      RECT 496.0500 0.0000 499.7500 0.6200 ;
      RECT 492.0500 0.0000 495.7500 0.6200 ;
      RECT 488.0500 0.0000 491.7500 0.6200 ;
      RECT 484.0500 0.0000 487.7500 0.6200 ;
      RECT 0.0000 0.0000 483.7500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 651.9500 1220.0000 1220.0000 ;
      RECT 0.6200 651.6500 1220.0000 651.9500 ;
      RECT 0.0000 647.9500 1220.0000 651.6500 ;
      RECT 0.6200 647.6500 1220.0000 647.9500 ;
      RECT 0.0000 643.9500 1220.0000 647.6500 ;
      RECT 0.6200 643.6500 1220.0000 643.9500 ;
      RECT 0.0000 639.9500 1220.0000 643.6500 ;
      RECT 0.6200 639.6500 1220.0000 639.9500 ;
      RECT 0.0000 635.9500 1220.0000 639.6500 ;
      RECT 0.6200 635.6500 1220.0000 635.9500 ;
      RECT 0.0000 631.9500 1220.0000 635.6500 ;
      RECT 0.6200 631.6500 1220.0000 631.9500 ;
      RECT 0.0000 627.9500 1220.0000 631.6500 ;
      RECT 0.6200 627.6500 1220.0000 627.9500 ;
      RECT 0.0000 623.9500 1220.0000 627.6500 ;
      RECT 0.6200 623.6500 1220.0000 623.9500 ;
      RECT 0.0000 619.9500 1220.0000 623.6500 ;
      RECT 0.6200 619.6500 1220.0000 619.9500 ;
      RECT 0.0000 615.9500 1220.0000 619.6500 ;
      RECT 0.6200 615.6500 1220.0000 615.9500 ;
      RECT 0.0000 611.9500 1220.0000 615.6500 ;
      RECT 0.6200 611.6500 1220.0000 611.9500 ;
      RECT 0.0000 607.9500 1220.0000 611.6500 ;
      RECT 0.6200 607.6500 1220.0000 607.9500 ;
      RECT 0.0000 603.9500 1220.0000 607.6500 ;
      RECT 0.6200 603.6500 1220.0000 603.9500 ;
      RECT 0.0000 599.9500 1220.0000 603.6500 ;
      RECT 0.6200 599.6500 1220.0000 599.9500 ;
      RECT 0.0000 595.9500 1220.0000 599.6500 ;
      RECT 0.6200 595.6500 1220.0000 595.9500 ;
      RECT 0.0000 591.9500 1220.0000 595.6500 ;
      RECT 0.6200 591.6500 1220.0000 591.9500 ;
      RECT 0.0000 587.9500 1220.0000 591.6500 ;
      RECT 0.6200 587.6500 1220.0000 587.9500 ;
      RECT 0.0000 583.9500 1220.0000 587.6500 ;
      RECT 0.6200 583.6500 1220.0000 583.9500 ;
      RECT 0.0000 579.9500 1220.0000 583.6500 ;
      RECT 0.6200 579.6500 1220.0000 579.9500 ;
      RECT 0.0000 575.9500 1220.0000 579.6500 ;
      RECT 0.6200 575.6500 1220.0000 575.9500 ;
      RECT 0.0000 571.9500 1220.0000 575.6500 ;
      RECT 0.6200 571.6500 1220.0000 571.9500 ;
      RECT 0.0000 567.9500 1220.0000 571.6500 ;
      RECT 0.6200 567.6500 1220.0000 567.9500 ;
      RECT 0.0000 0.0000 1220.0000 567.6500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 1220.0000 1220.0000 ;
    LAYER M5 ;
      RECT 0.0000 1210.2450 1220.0000 1220.0000 ;
      RECT 1214.5000 1207.2450 1220.0000 1210.2450 ;
      RECT 0.0000 1207.2450 5.5000 1210.2450 ;
      RECT 0.0000 1205.2450 1220.0000 1207.2450 ;
      RECT 1218.5000 1202.2450 1220.0000 1205.2450 ;
      RECT 0.0000 1202.2450 1.5000 1205.2450 ;
      RECT 0.0000 1202.2400 1220.0000 1202.2450 ;
      RECT 1214.5000 1199.2400 1220.0000 1202.2400 ;
      RECT 0.0000 1199.2400 5.5000 1202.2400 ;
      RECT 0.0000 1197.2400 1220.0000 1199.2400 ;
      RECT 1218.5000 1194.2400 1220.0000 1197.2400 ;
      RECT 0.0000 1194.2400 1.5000 1197.2400 ;
      RECT 0.0000 1194.2350 1220.0000 1194.2400 ;
      RECT 1214.5000 1191.2350 1220.0000 1194.2350 ;
      RECT 0.0000 1191.2350 5.5000 1194.2350 ;
      RECT 0.0000 1189.2350 1220.0000 1191.2350 ;
      RECT 1218.5000 1186.2350 1220.0000 1189.2350 ;
      RECT 0.0000 1186.2350 1.5000 1189.2350 ;
      RECT 0.0000 1186.2300 1220.0000 1186.2350 ;
      RECT 1214.5000 1183.2300 1220.0000 1186.2300 ;
      RECT 0.0000 1183.2300 5.5000 1186.2300 ;
      RECT 0.0000 1181.2300 1220.0000 1183.2300 ;
      RECT 1218.5000 1178.2300 1220.0000 1181.2300 ;
      RECT 0.0000 1178.2300 1.5000 1181.2300 ;
      RECT 0.0000 1178.2250 1220.0000 1178.2300 ;
      RECT 1214.5000 1175.2250 1220.0000 1178.2250 ;
      RECT 0.0000 1175.2250 5.5000 1178.2250 ;
      RECT 0.0000 1173.2250 1220.0000 1175.2250 ;
      RECT 1218.5000 1170.2250 1220.0000 1173.2250 ;
      RECT 0.0000 1170.2250 1.5000 1173.2250 ;
      RECT 0.0000 1170.2200 1220.0000 1170.2250 ;
      RECT 1214.5000 1167.2200 1220.0000 1170.2200 ;
      RECT 0.0000 1167.2200 5.5000 1170.2200 ;
      RECT 0.0000 1165.2200 1220.0000 1167.2200 ;
      RECT 1218.5000 1162.2200 1220.0000 1165.2200 ;
      RECT 0.0000 1162.2200 1.5000 1165.2200 ;
      RECT 0.0000 1162.2150 1220.0000 1162.2200 ;
      RECT 1214.5000 1159.2150 1220.0000 1162.2150 ;
      RECT 0.0000 1159.2150 5.5000 1162.2150 ;
      RECT 0.0000 1157.2150 1220.0000 1159.2150 ;
      RECT 1218.5000 1154.2150 1220.0000 1157.2150 ;
      RECT 0.0000 1154.2150 1.5000 1157.2150 ;
      RECT 0.0000 1154.2100 1220.0000 1154.2150 ;
      RECT 1214.5000 1151.2100 1220.0000 1154.2100 ;
      RECT 0.0000 1151.2100 5.5000 1154.2100 ;
      RECT 0.0000 1149.2100 1220.0000 1151.2100 ;
      RECT 1218.5000 1146.2100 1220.0000 1149.2100 ;
      RECT 0.0000 1146.2100 1.5000 1149.2100 ;
      RECT 0.0000 1146.2050 1220.0000 1146.2100 ;
      RECT 1214.5000 1143.2050 1220.0000 1146.2050 ;
      RECT 0.0000 1143.2050 5.5000 1146.2050 ;
      RECT 0.0000 1141.2050 1220.0000 1143.2050 ;
      RECT 1218.5000 1138.2050 1220.0000 1141.2050 ;
      RECT 0.0000 1138.2050 1.5000 1141.2050 ;
      RECT 0.0000 1138.2000 1220.0000 1138.2050 ;
      RECT 1214.5000 1135.2000 1220.0000 1138.2000 ;
      RECT 0.0000 1135.2000 5.5000 1138.2000 ;
      RECT 0.0000 1133.2000 1220.0000 1135.2000 ;
      RECT 1218.5000 1130.2000 1220.0000 1133.2000 ;
      RECT 0.0000 1130.2000 1.5000 1133.2000 ;
      RECT 0.0000 1130.1950 1220.0000 1130.2000 ;
      RECT 1214.5000 1127.1950 1220.0000 1130.1950 ;
      RECT 0.0000 1127.1950 5.5000 1130.1950 ;
      RECT 0.0000 1125.1950 1220.0000 1127.1950 ;
      RECT 1218.5000 1122.1950 1220.0000 1125.1950 ;
      RECT 0.0000 1122.1950 1.5000 1125.1950 ;
      RECT 0.0000 1122.1900 1220.0000 1122.1950 ;
      RECT 1214.5000 1119.1900 1220.0000 1122.1900 ;
      RECT 0.0000 1119.1900 5.5000 1122.1900 ;
      RECT 0.0000 1117.1900 1220.0000 1119.1900 ;
      RECT 1218.5000 1114.1900 1220.0000 1117.1900 ;
      RECT 0.0000 1114.1900 1.5000 1117.1900 ;
      RECT 0.0000 1114.1850 1220.0000 1114.1900 ;
      RECT 1214.5000 1111.1850 1220.0000 1114.1850 ;
      RECT 0.0000 1111.1850 5.5000 1114.1850 ;
      RECT 0.0000 1109.1850 1220.0000 1111.1850 ;
      RECT 1218.5000 1106.1850 1220.0000 1109.1850 ;
      RECT 0.0000 1106.1850 1.5000 1109.1850 ;
      RECT 0.0000 1106.1800 1220.0000 1106.1850 ;
      RECT 1214.5000 1103.1800 1220.0000 1106.1800 ;
      RECT 0.0000 1103.1800 5.5000 1106.1800 ;
      RECT 0.0000 1101.1800 1220.0000 1103.1800 ;
      RECT 1218.5000 1098.1800 1220.0000 1101.1800 ;
      RECT 0.0000 1098.1800 1.5000 1101.1800 ;
      RECT 0.0000 1098.1750 1220.0000 1098.1800 ;
      RECT 1214.5000 1095.1750 1220.0000 1098.1750 ;
      RECT 0.0000 1095.1750 5.5000 1098.1750 ;
      RECT 0.0000 1093.1750 1220.0000 1095.1750 ;
      RECT 1218.5000 1090.1750 1220.0000 1093.1750 ;
      RECT 0.0000 1090.1750 1.5000 1093.1750 ;
      RECT 0.0000 1090.1700 1220.0000 1090.1750 ;
      RECT 1214.5000 1087.1700 1220.0000 1090.1700 ;
      RECT 0.0000 1087.1700 5.5000 1090.1700 ;
      RECT 0.0000 1085.1700 1220.0000 1087.1700 ;
      RECT 1218.5000 1082.1700 1220.0000 1085.1700 ;
      RECT 0.0000 1082.1700 1.5000 1085.1700 ;
      RECT 0.0000 1082.1650 1220.0000 1082.1700 ;
      RECT 1214.5000 1079.1650 1220.0000 1082.1650 ;
      RECT 0.0000 1079.1650 5.5000 1082.1650 ;
      RECT 0.0000 1077.1650 1220.0000 1079.1650 ;
      RECT 1218.5000 1074.1650 1220.0000 1077.1650 ;
      RECT 0.0000 1074.1650 1.5000 1077.1650 ;
      RECT 0.0000 1074.1600 1220.0000 1074.1650 ;
      RECT 1214.5000 1071.1600 1220.0000 1074.1600 ;
      RECT 0.0000 1071.1600 5.5000 1074.1600 ;
      RECT 0.0000 1069.1600 1220.0000 1071.1600 ;
      RECT 1218.5000 1066.1600 1220.0000 1069.1600 ;
      RECT 0.0000 1066.1600 1.5000 1069.1600 ;
      RECT 0.0000 1066.1550 1220.0000 1066.1600 ;
      RECT 1214.5000 1063.1550 1220.0000 1066.1550 ;
      RECT 0.0000 1063.1550 5.5000 1066.1550 ;
      RECT 0.0000 1061.1550 1220.0000 1063.1550 ;
      RECT 1218.5000 1058.1550 1220.0000 1061.1550 ;
      RECT 0.0000 1058.1550 1.5000 1061.1550 ;
      RECT 0.0000 1058.1500 1220.0000 1058.1550 ;
      RECT 1214.5000 1055.1500 1220.0000 1058.1500 ;
      RECT 0.0000 1055.1500 5.5000 1058.1500 ;
      RECT 0.0000 1053.1500 1220.0000 1055.1500 ;
      RECT 1218.5000 1050.1500 1220.0000 1053.1500 ;
      RECT 0.0000 1050.1500 1.5000 1053.1500 ;
      RECT 0.0000 1050.1450 1220.0000 1050.1500 ;
      RECT 1214.5000 1047.1450 1220.0000 1050.1450 ;
      RECT 0.0000 1047.1450 5.5000 1050.1450 ;
      RECT 0.0000 1045.1450 1220.0000 1047.1450 ;
      RECT 1218.5000 1042.1450 1220.0000 1045.1450 ;
      RECT 0.0000 1042.1450 1.5000 1045.1450 ;
      RECT 0.0000 1042.1400 1220.0000 1042.1450 ;
      RECT 1214.5000 1039.1400 1220.0000 1042.1400 ;
      RECT 0.0000 1039.1400 5.5000 1042.1400 ;
      RECT 0.0000 1037.1400 1220.0000 1039.1400 ;
      RECT 1218.5000 1034.1400 1220.0000 1037.1400 ;
      RECT 0.0000 1034.1400 1.5000 1037.1400 ;
      RECT 0.0000 1034.1350 1220.0000 1034.1400 ;
      RECT 1214.5000 1031.1350 1220.0000 1034.1350 ;
      RECT 0.0000 1031.1350 5.5000 1034.1350 ;
      RECT 0.0000 1029.1350 1220.0000 1031.1350 ;
      RECT 1218.5000 1026.1350 1220.0000 1029.1350 ;
      RECT 0.0000 1026.1350 1.5000 1029.1350 ;
      RECT 0.0000 1026.1300 1220.0000 1026.1350 ;
      RECT 1214.5000 1023.1300 1220.0000 1026.1300 ;
      RECT 0.0000 1023.1300 5.5000 1026.1300 ;
      RECT 0.0000 1021.1300 1220.0000 1023.1300 ;
      RECT 1218.5000 1018.1300 1220.0000 1021.1300 ;
      RECT 0.0000 1018.1300 1.5000 1021.1300 ;
      RECT 0.0000 1018.1250 1220.0000 1018.1300 ;
      RECT 1214.5000 1015.1250 1220.0000 1018.1250 ;
      RECT 0.0000 1015.1250 5.5000 1018.1250 ;
      RECT 0.0000 1013.1250 1220.0000 1015.1250 ;
      RECT 1218.5000 1010.1250 1220.0000 1013.1250 ;
      RECT 0.0000 1010.1250 1.5000 1013.1250 ;
      RECT 0.0000 1010.1200 1220.0000 1010.1250 ;
      RECT 1214.5000 1007.1200 1220.0000 1010.1200 ;
      RECT 0.0000 1007.1200 5.5000 1010.1200 ;
      RECT 0.0000 1005.1200 1220.0000 1007.1200 ;
      RECT 1218.5000 1002.1200 1220.0000 1005.1200 ;
      RECT 0.0000 1002.1200 1.5000 1005.1200 ;
      RECT 0.0000 1002.1150 1220.0000 1002.1200 ;
      RECT 1214.5000 999.1150 1220.0000 1002.1150 ;
      RECT 0.0000 999.1150 5.5000 1002.1150 ;
      RECT 0.0000 997.1150 1220.0000 999.1150 ;
      RECT 1218.5000 994.1150 1220.0000 997.1150 ;
      RECT 0.0000 994.1150 1.5000 997.1150 ;
      RECT 0.0000 994.1100 1220.0000 994.1150 ;
      RECT 1214.5000 991.1100 1220.0000 994.1100 ;
      RECT 0.0000 991.1100 5.5000 994.1100 ;
      RECT 0.0000 989.1100 1220.0000 991.1100 ;
      RECT 1218.5000 986.1100 1220.0000 989.1100 ;
      RECT 0.0000 986.1100 1.5000 989.1100 ;
      RECT 0.0000 986.1050 1220.0000 986.1100 ;
      RECT 1214.5000 983.1050 1220.0000 986.1050 ;
      RECT 0.0000 983.1050 5.5000 986.1050 ;
      RECT 0.0000 981.1050 1220.0000 983.1050 ;
      RECT 1218.5000 978.1050 1220.0000 981.1050 ;
      RECT 0.0000 978.1050 1.5000 981.1050 ;
      RECT 0.0000 978.1000 1220.0000 978.1050 ;
      RECT 1214.5000 975.1000 1220.0000 978.1000 ;
      RECT 0.0000 975.1000 5.5000 978.1000 ;
      RECT 0.0000 973.1000 1220.0000 975.1000 ;
      RECT 1218.5000 970.1000 1220.0000 973.1000 ;
      RECT 0.0000 970.1000 1.5000 973.1000 ;
      RECT 0.0000 970.0950 1220.0000 970.1000 ;
      RECT 1214.5000 967.0950 1220.0000 970.0950 ;
      RECT 0.0000 967.0950 5.5000 970.0950 ;
      RECT 0.0000 965.0950 1220.0000 967.0950 ;
      RECT 1218.5000 962.0950 1220.0000 965.0950 ;
      RECT 0.0000 962.0950 1.5000 965.0950 ;
      RECT 0.0000 962.0900 1220.0000 962.0950 ;
      RECT 1214.5000 959.0900 1220.0000 962.0900 ;
      RECT 0.0000 959.0900 5.5000 962.0900 ;
      RECT 0.0000 957.0900 1220.0000 959.0900 ;
      RECT 1218.5000 954.0900 1220.0000 957.0900 ;
      RECT 0.0000 954.0900 1.5000 957.0900 ;
      RECT 0.0000 954.0850 1220.0000 954.0900 ;
      RECT 1214.5000 951.0850 1220.0000 954.0850 ;
      RECT 0.0000 951.0850 5.5000 954.0850 ;
      RECT 0.0000 949.0850 1220.0000 951.0850 ;
      RECT 1218.5000 946.0850 1220.0000 949.0850 ;
      RECT 0.0000 946.0850 1.5000 949.0850 ;
      RECT 0.0000 946.0800 1220.0000 946.0850 ;
      RECT 1214.5000 943.0800 1220.0000 946.0800 ;
      RECT 0.0000 943.0800 5.5000 946.0800 ;
      RECT 0.0000 941.0800 1220.0000 943.0800 ;
      RECT 1218.5000 938.0800 1220.0000 941.0800 ;
      RECT 0.0000 938.0800 1.5000 941.0800 ;
      RECT 0.0000 938.0750 1220.0000 938.0800 ;
      RECT 1214.5000 935.0750 1220.0000 938.0750 ;
      RECT 0.0000 935.0750 5.5000 938.0750 ;
      RECT 0.0000 933.0750 1220.0000 935.0750 ;
      RECT 1218.5000 930.0750 1220.0000 933.0750 ;
      RECT 0.0000 930.0750 1.5000 933.0750 ;
      RECT 0.0000 930.0700 1220.0000 930.0750 ;
      RECT 1214.5000 927.0700 1220.0000 930.0700 ;
      RECT 0.0000 927.0700 5.5000 930.0700 ;
      RECT 0.0000 925.0700 1220.0000 927.0700 ;
      RECT 1218.5000 922.0700 1220.0000 925.0700 ;
      RECT 0.0000 922.0700 1.5000 925.0700 ;
      RECT 0.0000 922.0650 1220.0000 922.0700 ;
      RECT 1214.5000 919.0650 1220.0000 922.0650 ;
      RECT 0.0000 919.0650 5.5000 922.0650 ;
      RECT 0.0000 917.0650 1220.0000 919.0650 ;
      RECT 1218.5000 914.0650 1220.0000 917.0650 ;
      RECT 0.0000 914.0650 1.5000 917.0650 ;
      RECT 0.0000 914.0600 1220.0000 914.0650 ;
      RECT 1214.5000 911.0600 1220.0000 914.0600 ;
      RECT 0.0000 911.0600 5.5000 914.0600 ;
      RECT 0.0000 909.0600 1220.0000 911.0600 ;
      RECT 1218.5000 906.0600 1220.0000 909.0600 ;
      RECT 0.0000 906.0600 1.5000 909.0600 ;
      RECT 0.0000 906.0550 1220.0000 906.0600 ;
      RECT 1214.5000 903.0550 1220.0000 906.0550 ;
      RECT 0.0000 903.0550 5.5000 906.0550 ;
      RECT 0.0000 901.0550 1220.0000 903.0550 ;
      RECT 1218.5000 898.0550 1220.0000 901.0550 ;
      RECT 0.0000 898.0550 1.5000 901.0550 ;
      RECT 0.0000 898.0500 1220.0000 898.0550 ;
      RECT 1214.5000 895.0500 1220.0000 898.0500 ;
      RECT 0.0000 895.0500 5.5000 898.0500 ;
      RECT 0.0000 893.0500 1220.0000 895.0500 ;
      RECT 1218.5000 890.0500 1220.0000 893.0500 ;
      RECT 0.0000 890.0500 1.5000 893.0500 ;
      RECT 0.0000 890.0450 1220.0000 890.0500 ;
      RECT 1214.5000 887.0450 1220.0000 890.0450 ;
      RECT 0.0000 887.0450 5.5000 890.0450 ;
      RECT 0.0000 885.0450 1220.0000 887.0450 ;
      RECT 1218.5000 882.0450 1220.0000 885.0450 ;
      RECT 0.0000 882.0450 1.5000 885.0450 ;
      RECT 0.0000 882.0400 1220.0000 882.0450 ;
      RECT 1214.5000 879.0400 1220.0000 882.0400 ;
      RECT 0.0000 879.0400 5.5000 882.0400 ;
      RECT 0.0000 877.0400 1220.0000 879.0400 ;
      RECT 1218.5000 874.0400 1220.0000 877.0400 ;
      RECT 0.0000 874.0400 1.5000 877.0400 ;
      RECT 0.0000 874.0350 1220.0000 874.0400 ;
      RECT 1214.5000 871.0350 1220.0000 874.0350 ;
      RECT 0.0000 871.0350 5.5000 874.0350 ;
      RECT 0.0000 869.0350 1220.0000 871.0350 ;
      RECT 1218.5000 866.0350 1220.0000 869.0350 ;
      RECT 0.0000 866.0350 1.5000 869.0350 ;
      RECT 0.0000 866.0300 1220.0000 866.0350 ;
      RECT 1214.5000 863.0300 1220.0000 866.0300 ;
      RECT 0.0000 863.0300 5.5000 866.0300 ;
      RECT 0.0000 861.0300 1220.0000 863.0300 ;
      RECT 1218.5000 858.0300 1220.0000 861.0300 ;
      RECT 0.0000 858.0300 1.5000 861.0300 ;
      RECT 0.0000 858.0250 1220.0000 858.0300 ;
      RECT 1214.5000 855.0250 1220.0000 858.0250 ;
      RECT 0.0000 855.0250 5.5000 858.0250 ;
      RECT 0.0000 853.0250 1220.0000 855.0250 ;
      RECT 1218.5000 850.0250 1220.0000 853.0250 ;
      RECT 0.0000 850.0250 1.5000 853.0250 ;
      RECT 0.0000 850.0200 1220.0000 850.0250 ;
      RECT 1214.5000 847.0200 1220.0000 850.0200 ;
      RECT 0.0000 847.0200 5.5000 850.0200 ;
      RECT 0.0000 845.0200 1220.0000 847.0200 ;
      RECT 1218.5000 842.0200 1220.0000 845.0200 ;
      RECT 0.0000 842.0200 1.5000 845.0200 ;
      RECT 0.0000 842.0150 1220.0000 842.0200 ;
      RECT 1214.5000 839.0150 1220.0000 842.0150 ;
      RECT 0.0000 839.0150 5.5000 842.0150 ;
      RECT 0.0000 837.0150 1220.0000 839.0150 ;
      RECT 1218.5000 834.0150 1220.0000 837.0150 ;
      RECT 0.0000 834.0150 1.5000 837.0150 ;
      RECT 0.0000 834.0100 1220.0000 834.0150 ;
      RECT 1214.5000 831.0100 1220.0000 834.0100 ;
      RECT 0.0000 831.0100 5.5000 834.0100 ;
      RECT 0.0000 829.0100 1220.0000 831.0100 ;
      RECT 1218.5000 826.0100 1220.0000 829.0100 ;
      RECT 0.0000 826.0100 1.5000 829.0100 ;
      RECT 0.0000 826.0050 1220.0000 826.0100 ;
      RECT 1214.5000 823.0050 1220.0000 826.0050 ;
      RECT 0.0000 823.0050 5.5000 826.0050 ;
      RECT 0.0000 821.0050 1220.0000 823.0050 ;
      RECT 1218.5000 818.0050 1220.0000 821.0050 ;
      RECT 0.0000 818.0050 1.5000 821.0050 ;
      RECT 0.0000 818.0000 1220.0000 818.0050 ;
      RECT 1214.5000 815.0000 1220.0000 818.0000 ;
      RECT 0.0000 815.0000 5.5000 818.0000 ;
      RECT 0.0000 813.0000 1220.0000 815.0000 ;
      RECT 1218.5000 810.0000 1220.0000 813.0000 ;
      RECT 0.0000 810.0000 1.5000 813.0000 ;
      RECT 0.0000 809.9950 1220.0000 810.0000 ;
      RECT 1214.5000 806.9950 1220.0000 809.9950 ;
      RECT 0.0000 806.9950 5.5000 809.9950 ;
      RECT 0.0000 804.9950 1220.0000 806.9950 ;
      RECT 1218.5000 801.9950 1220.0000 804.9950 ;
      RECT 0.0000 801.9950 1.5000 804.9950 ;
      RECT 0.0000 801.9900 1220.0000 801.9950 ;
      RECT 1214.5000 798.9900 1220.0000 801.9900 ;
      RECT 0.0000 798.9900 5.5000 801.9900 ;
      RECT 0.0000 796.9900 1220.0000 798.9900 ;
      RECT 1218.5000 793.9900 1220.0000 796.9900 ;
      RECT 0.0000 793.9900 1.5000 796.9900 ;
      RECT 0.0000 793.9850 1220.0000 793.9900 ;
      RECT 1214.5000 790.9850 1220.0000 793.9850 ;
      RECT 0.0000 790.9850 5.5000 793.9850 ;
      RECT 0.0000 788.9850 1220.0000 790.9850 ;
      RECT 1218.5000 785.9850 1220.0000 788.9850 ;
      RECT 0.0000 785.9850 1.5000 788.9850 ;
      RECT 0.0000 785.9800 1220.0000 785.9850 ;
      RECT 1214.5000 782.9800 1220.0000 785.9800 ;
      RECT 0.0000 782.9800 5.5000 785.9800 ;
      RECT 0.0000 780.9800 1220.0000 782.9800 ;
      RECT 1218.5000 777.9800 1220.0000 780.9800 ;
      RECT 0.0000 777.9800 1.5000 780.9800 ;
      RECT 0.0000 777.9750 1220.0000 777.9800 ;
      RECT 1214.5000 774.9750 1220.0000 777.9750 ;
      RECT 0.0000 774.9750 5.5000 777.9750 ;
      RECT 0.0000 772.9750 1220.0000 774.9750 ;
      RECT 1218.5000 769.9750 1220.0000 772.9750 ;
      RECT 0.0000 769.9750 1.5000 772.9750 ;
      RECT 0.0000 769.9700 1220.0000 769.9750 ;
      RECT 1214.5000 766.9700 1220.0000 769.9700 ;
      RECT 0.0000 766.9700 5.5000 769.9700 ;
      RECT 0.0000 764.9700 1220.0000 766.9700 ;
      RECT 1218.5000 761.9700 1220.0000 764.9700 ;
      RECT 0.0000 761.9700 1.5000 764.9700 ;
      RECT 0.0000 761.9650 1220.0000 761.9700 ;
      RECT 1214.5000 758.9650 1220.0000 761.9650 ;
      RECT 0.0000 758.9650 5.5000 761.9650 ;
      RECT 0.0000 756.9650 1220.0000 758.9650 ;
      RECT 1218.5000 753.9650 1220.0000 756.9650 ;
      RECT 0.0000 753.9650 1.5000 756.9650 ;
      RECT 0.0000 753.9600 1220.0000 753.9650 ;
      RECT 1214.5000 750.9600 1220.0000 753.9600 ;
      RECT 0.0000 750.9600 5.5000 753.9600 ;
      RECT 0.0000 748.9600 1220.0000 750.9600 ;
      RECT 1218.5000 745.9600 1220.0000 748.9600 ;
      RECT 0.0000 745.9600 1.5000 748.9600 ;
      RECT 0.0000 745.9550 1220.0000 745.9600 ;
      RECT 1214.5000 742.9550 1220.0000 745.9550 ;
      RECT 0.0000 742.9550 5.5000 745.9550 ;
      RECT 0.0000 740.9550 1220.0000 742.9550 ;
      RECT 1218.5000 737.9550 1220.0000 740.9550 ;
      RECT 0.0000 737.9550 1.5000 740.9550 ;
      RECT 0.0000 737.9500 1220.0000 737.9550 ;
      RECT 1214.5000 734.9500 1220.0000 737.9500 ;
      RECT 0.0000 734.9500 5.5000 737.9500 ;
      RECT 0.0000 732.9500 1220.0000 734.9500 ;
      RECT 1218.5000 729.9500 1220.0000 732.9500 ;
      RECT 0.0000 729.9500 1.5000 732.9500 ;
      RECT 0.0000 729.9450 1220.0000 729.9500 ;
      RECT 1214.5000 726.9450 1220.0000 729.9450 ;
      RECT 0.0000 726.9450 5.5000 729.9450 ;
      RECT 0.0000 724.9450 1220.0000 726.9450 ;
      RECT 1218.5000 721.9450 1220.0000 724.9450 ;
      RECT 0.0000 721.9450 1.5000 724.9450 ;
      RECT 0.0000 721.9400 1220.0000 721.9450 ;
      RECT 1214.5000 718.9400 1220.0000 721.9400 ;
      RECT 0.0000 718.9400 5.5000 721.9400 ;
      RECT 0.0000 716.9400 1220.0000 718.9400 ;
      RECT 1218.5000 713.9400 1220.0000 716.9400 ;
      RECT 0.0000 713.9400 1.5000 716.9400 ;
      RECT 0.0000 713.9350 1220.0000 713.9400 ;
      RECT 1214.5000 710.9350 1220.0000 713.9350 ;
      RECT 0.0000 710.9350 5.5000 713.9350 ;
      RECT 0.0000 708.9350 1220.0000 710.9350 ;
      RECT 1218.5000 705.9350 1220.0000 708.9350 ;
      RECT 0.0000 705.9350 1.5000 708.9350 ;
      RECT 0.0000 705.9300 1220.0000 705.9350 ;
      RECT 1214.5000 702.9300 1220.0000 705.9300 ;
      RECT 0.0000 702.9300 5.5000 705.9300 ;
      RECT 0.0000 700.9300 1220.0000 702.9300 ;
      RECT 1218.5000 697.9300 1220.0000 700.9300 ;
      RECT 0.0000 697.9300 1.5000 700.9300 ;
      RECT 0.0000 697.9250 1220.0000 697.9300 ;
      RECT 1214.5000 694.9250 1220.0000 697.9250 ;
      RECT 0.0000 694.9250 5.5000 697.9250 ;
      RECT 0.0000 692.9250 1220.0000 694.9250 ;
      RECT 1218.5000 689.9250 1220.0000 692.9250 ;
      RECT 0.0000 689.9250 1.5000 692.9250 ;
      RECT 0.0000 689.9200 1220.0000 689.9250 ;
      RECT 1214.5000 686.9200 1220.0000 689.9200 ;
      RECT 0.0000 686.9200 5.5000 689.9200 ;
      RECT 0.0000 684.9200 1220.0000 686.9200 ;
      RECT 1218.5000 681.9200 1220.0000 684.9200 ;
      RECT 0.0000 681.9200 1.5000 684.9200 ;
      RECT 0.0000 681.9150 1220.0000 681.9200 ;
      RECT 1214.5000 678.9150 1220.0000 681.9150 ;
      RECT 0.0000 678.9150 5.5000 681.9150 ;
      RECT 0.0000 676.9150 1220.0000 678.9150 ;
      RECT 1218.5000 673.9150 1220.0000 676.9150 ;
      RECT 0.0000 673.9150 1.5000 676.9150 ;
      RECT 0.0000 673.9100 1220.0000 673.9150 ;
      RECT 1214.5000 670.9100 1220.0000 673.9100 ;
      RECT 0.0000 670.9100 5.5000 673.9100 ;
      RECT 0.0000 668.9100 1220.0000 670.9100 ;
      RECT 1218.5000 665.9100 1220.0000 668.9100 ;
      RECT 0.0000 665.9100 1.5000 668.9100 ;
      RECT 0.0000 665.9050 1220.0000 665.9100 ;
      RECT 1214.5000 662.9050 1220.0000 665.9050 ;
      RECT 0.0000 662.9050 5.5000 665.9050 ;
      RECT 0.0000 660.9050 1220.0000 662.9050 ;
      RECT 1218.5000 657.9050 1220.0000 660.9050 ;
      RECT 0.0000 657.9050 1.5000 660.9050 ;
      RECT 0.0000 657.9000 1220.0000 657.9050 ;
      RECT 1214.5000 654.9000 1220.0000 657.9000 ;
      RECT 0.0000 654.9000 5.5000 657.9000 ;
      RECT 0.0000 652.9000 1220.0000 654.9000 ;
      RECT 1218.5000 649.9000 1220.0000 652.9000 ;
      RECT 0.0000 649.9000 1.5000 652.9000 ;
      RECT 0.0000 649.8950 1220.0000 649.9000 ;
      RECT 1214.5000 646.8950 1220.0000 649.8950 ;
      RECT 0.0000 646.8950 5.5000 649.8950 ;
      RECT 0.0000 644.8950 1220.0000 646.8950 ;
      RECT 1218.5000 641.8950 1220.0000 644.8950 ;
      RECT 0.0000 641.8950 1.5000 644.8950 ;
      RECT 0.0000 641.8900 1220.0000 641.8950 ;
      RECT 1214.5000 638.8900 1220.0000 641.8900 ;
      RECT 0.0000 638.8900 5.5000 641.8900 ;
      RECT 0.0000 636.8900 1220.0000 638.8900 ;
      RECT 1218.5000 633.8900 1220.0000 636.8900 ;
      RECT 0.0000 633.8900 1.5000 636.8900 ;
      RECT 0.0000 633.8850 1220.0000 633.8900 ;
      RECT 1214.5000 630.8850 1220.0000 633.8850 ;
      RECT 0.0000 630.8850 5.5000 633.8850 ;
      RECT 0.0000 628.8850 1220.0000 630.8850 ;
      RECT 1218.5000 625.8850 1220.0000 628.8850 ;
      RECT 0.0000 625.8850 1.5000 628.8850 ;
      RECT 0.0000 625.8800 1220.0000 625.8850 ;
      RECT 1214.5000 622.8800 1220.0000 625.8800 ;
      RECT 0.0000 622.8800 5.5000 625.8800 ;
      RECT 0.0000 620.8800 1220.0000 622.8800 ;
      RECT 1218.5000 617.8800 1220.0000 620.8800 ;
      RECT 0.0000 617.8800 1.5000 620.8800 ;
      RECT 0.0000 617.8750 1220.0000 617.8800 ;
      RECT 1214.5000 614.8750 1220.0000 617.8750 ;
      RECT 0.0000 614.8750 5.5000 617.8750 ;
      RECT 0.0000 612.8750 1220.0000 614.8750 ;
      RECT 1218.5000 609.8750 1220.0000 612.8750 ;
      RECT 0.0000 609.8750 1.5000 612.8750 ;
      RECT 0.0000 609.8700 1220.0000 609.8750 ;
      RECT 1214.5000 606.8700 1220.0000 609.8700 ;
      RECT 0.0000 606.8700 5.5000 609.8700 ;
      RECT 0.0000 604.8700 1220.0000 606.8700 ;
      RECT 1218.5000 601.8700 1220.0000 604.8700 ;
      RECT 0.0000 601.8700 1.5000 604.8700 ;
      RECT 0.0000 601.8650 1220.0000 601.8700 ;
      RECT 1214.5000 598.8650 1220.0000 601.8650 ;
      RECT 0.0000 598.8650 5.5000 601.8650 ;
      RECT 0.0000 596.8650 1220.0000 598.8650 ;
      RECT 1218.5000 593.8650 1220.0000 596.8650 ;
      RECT 0.0000 593.8650 1.5000 596.8650 ;
      RECT 0.0000 593.8600 1220.0000 593.8650 ;
      RECT 1214.5000 590.8600 1220.0000 593.8600 ;
      RECT 0.0000 590.8600 5.5000 593.8600 ;
      RECT 0.0000 588.8600 1220.0000 590.8600 ;
      RECT 1218.5000 585.8600 1220.0000 588.8600 ;
      RECT 0.0000 585.8600 1.5000 588.8600 ;
      RECT 0.0000 585.8550 1220.0000 585.8600 ;
      RECT 1214.5000 582.8550 1220.0000 585.8550 ;
      RECT 0.0000 582.8550 5.5000 585.8550 ;
      RECT 0.0000 580.8550 1220.0000 582.8550 ;
      RECT 1218.5000 577.8550 1220.0000 580.8550 ;
      RECT 0.0000 577.8550 1.5000 580.8550 ;
      RECT 0.0000 577.8500 1220.0000 577.8550 ;
      RECT 1214.5000 574.8500 1220.0000 577.8500 ;
      RECT 0.0000 574.8500 5.5000 577.8500 ;
      RECT 0.0000 572.8500 1220.0000 574.8500 ;
      RECT 1218.5000 569.8500 1220.0000 572.8500 ;
      RECT 0.0000 569.8500 1.5000 572.8500 ;
      RECT 0.0000 569.8450 1220.0000 569.8500 ;
      RECT 1214.5000 566.8450 1220.0000 569.8450 ;
      RECT 0.0000 566.8450 5.5000 569.8450 ;
      RECT 0.0000 564.8450 1220.0000 566.8450 ;
      RECT 1218.5000 561.8450 1220.0000 564.8450 ;
      RECT 0.0000 561.8450 1.5000 564.8450 ;
      RECT 0.0000 561.8400 1220.0000 561.8450 ;
      RECT 1214.5000 558.8400 1220.0000 561.8400 ;
      RECT 0.0000 558.8400 5.5000 561.8400 ;
      RECT 0.0000 556.8400 1220.0000 558.8400 ;
      RECT 1218.5000 553.8400 1220.0000 556.8400 ;
      RECT 0.0000 553.8400 1.5000 556.8400 ;
      RECT 0.0000 553.8350 1220.0000 553.8400 ;
      RECT 1214.5000 550.8350 1220.0000 553.8350 ;
      RECT 0.0000 550.8350 5.5000 553.8350 ;
      RECT 0.0000 548.8350 1220.0000 550.8350 ;
      RECT 1218.5000 545.8350 1220.0000 548.8350 ;
      RECT 0.0000 545.8350 1.5000 548.8350 ;
      RECT 0.0000 545.8300 1220.0000 545.8350 ;
      RECT 1214.5000 542.8300 1220.0000 545.8300 ;
      RECT 0.0000 542.8300 5.5000 545.8300 ;
      RECT 0.0000 540.8300 1220.0000 542.8300 ;
      RECT 1218.5000 537.8300 1220.0000 540.8300 ;
      RECT 0.0000 537.8300 1.5000 540.8300 ;
      RECT 0.0000 537.8250 1220.0000 537.8300 ;
      RECT 1214.5000 534.8250 1220.0000 537.8250 ;
      RECT 0.0000 534.8250 5.5000 537.8250 ;
      RECT 0.0000 532.8250 1220.0000 534.8250 ;
      RECT 1218.5000 529.8250 1220.0000 532.8250 ;
      RECT 0.0000 529.8250 1.5000 532.8250 ;
      RECT 0.0000 529.8200 1220.0000 529.8250 ;
      RECT 1214.5000 526.8200 1220.0000 529.8200 ;
      RECT 0.0000 526.8200 5.5000 529.8200 ;
      RECT 0.0000 524.8200 1220.0000 526.8200 ;
      RECT 1218.5000 521.8200 1220.0000 524.8200 ;
      RECT 0.0000 521.8200 1.5000 524.8200 ;
      RECT 0.0000 521.8150 1220.0000 521.8200 ;
      RECT 1214.5000 518.8150 1220.0000 521.8150 ;
      RECT 0.0000 518.8150 5.5000 521.8150 ;
      RECT 0.0000 516.8150 1220.0000 518.8150 ;
      RECT 1218.5000 513.8150 1220.0000 516.8150 ;
      RECT 0.0000 513.8150 1.5000 516.8150 ;
      RECT 0.0000 513.8100 1220.0000 513.8150 ;
      RECT 1214.5000 510.8100 1220.0000 513.8100 ;
      RECT 0.0000 510.8100 5.5000 513.8100 ;
      RECT 0.0000 508.8100 1220.0000 510.8100 ;
      RECT 1218.5000 505.8100 1220.0000 508.8100 ;
      RECT 0.0000 505.8100 1.5000 508.8100 ;
      RECT 0.0000 505.8050 1220.0000 505.8100 ;
      RECT 1214.5000 502.8050 1220.0000 505.8050 ;
      RECT 0.0000 502.8050 5.5000 505.8050 ;
      RECT 0.0000 500.8050 1220.0000 502.8050 ;
      RECT 1218.5000 497.8050 1220.0000 500.8050 ;
      RECT 0.0000 497.8050 1.5000 500.8050 ;
      RECT 0.0000 497.8000 1220.0000 497.8050 ;
      RECT 1214.5000 494.8000 1220.0000 497.8000 ;
      RECT 0.0000 494.8000 5.5000 497.8000 ;
      RECT 0.0000 492.8000 1220.0000 494.8000 ;
      RECT 1218.5000 489.8000 1220.0000 492.8000 ;
      RECT 0.0000 489.8000 1.5000 492.8000 ;
      RECT 0.0000 489.7950 1220.0000 489.8000 ;
      RECT 1214.5000 486.7950 1220.0000 489.7950 ;
      RECT 0.0000 486.7950 5.5000 489.7950 ;
      RECT 0.0000 484.7950 1220.0000 486.7950 ;
      RECT 1218.5000 481.7950 1220.0000 484.7950 ;
      RECT 0.0000 481.7950 1.5000 484.7950 ;
      RECT 0.0000 481.7900 1220.0000 481.7950 ;
      RECT 1214.5000 478.7900 1220.0000 481.7900 ;
      RECT 0.0000 478.7900 5.5000 481.7900 ;
      RECT 0.0000 476.7900 1220.0000 478.7900 ;
      RECT 1218.5000 473.7900 1220.0000 476.7900 ;
      RECT 0.0000 473.7900 1.5000 476.7900 ;
      RECT 0.0000 473.7850 1220.0000 473.7900 ;
      RECT 1214.5000 470.7850 1220.0000 473.7850 ;
      RECT 0.0000 470.7850 5.5000 473.7850 ;
      RECT 0.0000 468.7850 1220.0000 470.7850 ;
      RECT 1218.5000 465.7850 1220.0000 468.7850 ;
      RECT 0.0000 465.7850 1.5000 468.7850 ;
      RECT 0.0000 465.7800 1220.0000 465.7850 ;
      RECT 1214.5000 462.7800 1220.0000 465.7800 ;
      RECT 0.0000 462.7800 5.5000 465.7800 ;
      RECT 0.0000 460.7800 1220.0000 462.7800 ;
      RECT 1218.5000 457.7800 1220.0000 460.7800 ;
      RECT 0.0000 457.7800 1.5000 460.7800 ;
      RECT 0.0000 457.7750 1220.0000 457.7800 ;
      RECT 1214.5000 454.7750 1220.0000 457.7750 ;
      RECT 0.0000 454.7750 5.5000 457.7750 ;
      RECT 0.0000 452.7750 1220.0000 454.7750 ;
      RECT 1218.5000 449.7750 1220.0000 452.7750 ;
      RECT 0.0000 449.7750 1.5000 452.7750 ;
      RECT 0.0000 449.7700 1220.0000 449.7750 ;
      RECT 1214.5000 446.7700 1220.0000 449.7700 ;
      RECT 0.0000 446.7700 5.5000 449.7700 ;
      RECT 0.0000 444.7700 1220.0000 446.7700 ;
      RECT 1218.5000 441.7700 1220.0000 444.7700 ;
      RECT 0.0000 441.7700 1.5000 444.7700 ;
      RECT 0.0000 441.7650 1220.0000 441.7700 ;
      RECT 1214.5000 438.7650 1220.0000 441.7650 ;
      RECT 0.0000 438.7650 5.5000 441.7650 ;
      RECT 0.0000 436.7650 1220.0000 438.7650 ;
      RECT 1218.5000 433.7650 1220.0000 436.7650 ;
      RECT 0.0000 433.7650 1.5000 436.7650 ;
      RECT 0.0000 433.7600 1220.0000 433.7650 ;
      RECT 1214.5000 430.7600 1220.0000 433.7600 ;
      RECT 0.0000 430.7600 5.5000 433.7600 ;
      RECT 0.0000 428.7600 1220.0000 430.7600 ;
      RECT 1218.5000 425.7600 1220.0000 428.7600 ;
      RECT 0.0000 425.7600 1.5000 428.7600 ;
      RECT 0.0000 425.7550 1220.0000 425.7600 ;
      RECT 1214.5000 422.7550 1220.0000 425.7550 ;
      RECT 0.0000 422.7550 5.5000 425.7550 ;
      RECT 0.0000 420.7550 1220.0000 422.7550 ;
      RECT 1218.5000 417.7550 1220.0000 420.7550 ;
      RECT 0.0000 417.7550 1.5000 420.7550 ;
      RECT 0.0000 417.7500 1220.0000 417.7550 ;
      RECT 1214.5000 414.7500 1220.0000 417.7500 ;
      RECT 0.0000 414.7500 5.5000 417.7500 ;
      RECT 0.0000 412.7500 1220.0000 414.7500 ;
      RECT 1218.5000 409.7500 1220.0000 412.7500 ;
      RECT 0.0000 409.7500 1.5000 412.7500 ;
      RECT 0.0000 409.7450 1220.0000 409.7500 ;
      RECT 1214.5000 406.7450 1220.0000 409.7450 ;
      RECT 0.0000 406.7450 5.5000 409.7450 ;
      RECT 0.0000 404.7450 1220.0000 406.7450 ;
      RECT 1218.5000 401.7450 1220.0000 404.7450 ;
      RECT 0.0000 401.7450 1.5000 404.7450 ;
      RECT 0.0000 401.7400 1220.0000 401.7450 ;
      RECT 1214.5000 398.7400 1220.0000 401.7400 ;
      RECT 0.0000 398.7400 5.5000 401.7400 ;
      RECT 0.0000 396.7400 1220.0000 398.7400 ;
      RECT 1218.5000 393.7400 1220.0000 396.7400 ;
      RECT 0.0000 393.7400 1.5000 396.7400 ;
      RECT 0.0000 393.7350 1220.0000 393.7400 ;
      RECT 1214.5000 390.7350 1220.0000 393.7350 ;
      RECT 0.0000 390.7350 5.5000 393.7350 ;
      RECT 0.0000 388.7350 1220.0000 390.7350 ;
      RECT 1218.5000 385.7350 1220.0000 388.7350 ;
      RECT 0.0000 385.7350 1.5000 388.7350 ;
      RECT 0.0000 385.7300 1220.0000 385.7350 ;
      RECT 1214.5000 382.7300 1220.0000 385.7300 ;
      RECT 0.0000 382.7300 5.5000 385.7300 ;
      RECT 0.0000 380.7300 1220.0000 382.7300 ;
      RECT 1218.5000 377.7300 1220.0000 380.7300 ;
      RECT 0.0000 377.7300 1.5000 380.7300 ;
      RECT 0.0000 377.7250 1220.0000 377.7300 ;
      RECT 1214.5000 374.7250 1220.0000 377.7250 ;
      RECT 0.0000 374.7250 5.5000 377.7250 ;
      RECT 0.0000 372.7250 1220.0000 374.7250 ;
      RECT 1218.5000 369.7250 1220.0000 372.7250 ;
      RECT 0.0000 369.7250 1.5000 372.7250 ;
      RECT 0.0000 369.7200 1220.0000 369.7250 ;
      RECT 1214.5000 366.7200 1220.0000 369.7200 ;
      RECT 0.0000 366.7200 5.5000 369.7200 ;
      RECT 0.0000 364.7200 1220.0000 366.7200 ;
      RECT 1218.5000 361.7200 1220.0000 364.7200 ;
      RECT 0.0000 361.7200 1.5000 364.7200 ;
      RECT 0.0000 361.7150 1220.0000 361.7200 ;
      RECT 1214.5000 358.7150 1220.0000 361.7150 ;
      RECT 0.0000 358.7150 5.5000 361.7150 ;
      RECT 0.0000 356.7150 1220.0000 358.7150 ;
      RECT 1218.5000 353.7150 1220.0000 356.7150 ;
      RECT 0.0000 353.7150 1.5000 356.7150 ;
      RECT 0.0000 353.7100 1220.0000 353.7150 ;
      RECT 1214.5000 350.7100 1220.0000 353.7100 ;
      RECT 0.0000 350.7100 5.5000 353.7100 ;
      RECT 0.0000 348.7100 1220.0000 350.7100 ;
      RECT 1218.5000 345.7100 1220.0000 348.7100 ;
      RECT 0.0000 345.7100 1.5000 348.7100 ;
      RECT 0.0000 345.7050 1220.0000 345.7100 ;
      RECT 1214.5000 342.7050 1220.0000 345.7050 ;
      RECT 0.0000 342.7050 5.5000 345.7050 ;
      RECT 0.0000 340.7050 1220.0000 342.7050 ;
      RECT 1218.5000 337.7050 1220.0000 340.7050 ;
      RECT 0.0000 337.7050 1.5000 340.7050 ;
      RECT 0.0000 337.7000 1220.0000 337.7050 ;
      RECT 1214.5000 334.7000 1220.0000 337.7000 ;
      RECT 0.0000 334.7000 5.5000 337.7000 ;
      RECT 0.0000 332.7000 1220.0000 334.7000 ;
      RECT 1218.5000 329.7000 1220.0000 332.7000 ;
      RECT 0.0000 329.7000 1.5000 332.7000 ;
      RECT 0.0000 329.6950 1220.0000 329.7000 ;
      RECT 1214.5000 326.6950 1220.0000 329.6950 ;
      RECT 0.0000 326.6950 5.5000 329.6950 ;
      RECT 0.0000 324.6950 1220.0000 326.6950 ;
      RECT 1218.5000 321.6950 1220.0000 324.6950 ;
      RECT 0.0000 321.6950 1.5000 324.6950 ;
      RECT 0.0000 321.6900 1220.0000 321.6950 ;
      RECT 1214.5000 318.6900 1220.0000 321.6900 ;
      RECT 0.0000 318.6900 5.5000 321.6900 ;
      RECT 0.0000 316.6900 1220.0000 318.6900 ;
      RECT 1218.5000 313.6900 1220.0000 316.6900 ;
      RECT 0.0000 313.6900 1.5000 316.6900 ;
      RECT 0.0000 313.6850 1220.0000 313.6900 ;
      RECT 1214.5000 310.6850 1220.0000 313.6850 ;
      RECT 0.0000 310.6850 5.5000 313.6850 ;
      RECT 0.0000 308.6850 1220.0000 310.6850 ;
      RECT 1218.5000 305.6850 1220.0000 308.6850 ;
      RECT 0.0000 305.6850 1.5000 308.6850 ;
      RECT 0.0000 305.6800 1220.0000 305.6850 ;
      RECT 1214.5000 302.6800 1220.0000 305.6800 ;
      RECT 0.0000 302.6800 5.5000 305.6800 ;
      RECT 0.0000 300.6800 1220.0000 302.6800 ;
      RECT 1218.5000 297.6800 1220.0000 300.6800 ;
      RECT 0.0000 297.6800 1.5000 300.6800 ;
      RECT 0.0000 297.6750 1220.0000 297.6800 ;
      RECT 1214.5000 294.6750 1220.0000 297.6750 ;
      RECT 0.0000 294.6750 5.5000 297.6750 ;
      RECT 0.0000 292.6750 1220.0000 294.6750 ;
      RECT 1218.5000 289.6750 1220.0000 292.6750 ;
      RECT 0.0000 289.6750 1.5000 292.6750 ;
      RECT 0.0000 289.6700 1220.0000 289.6750 ;
      RECT 1214.5000 286.6700 1220.0000 289.6700 ;
      RECT 0.0000 286.6700 5.5000 289.6700 ;
      RECT 0.0000 284.6700 1220.0000 286.6700 ;
      RECT 1218.5000 281.6700 1220.0000 284.6700 ;
      RECT 0.0000 281.6700 1.5000 284.6700 ;
      RECT 0.0000 281.6650 1220.0000 281.6700 ;
      RECT 1214.5000 278.6650 1220.0000 281.6650 ;
      RECT 0.0000 278.6650 5.5000 281.6650 ;
      RECT 0.0000 276.6650 1220.0000 278.6650 ;
      RECT 1218.5000 273.6650 1220.0000 276.6650 ;
      RECT 0.0000 273.6650 1.5000 276.6650 ;
      RECT 0.0000 273.6600 1220.0000 273.6650 ;
      RECT 1214.5000 270.6600 1220.0000 273.6600 ;
      RECT 0.0000 270.6600 5.5000 273.6600 ;
      RECT 0.0000 268.6600 1220.0000 270.6600 ;
      RECT 1218.5000 265.6600 1220.0000 268.6600 ;
      RECT 0.0000 265.6600 1.5000 268.6600 ;
      RECT 0.0000 265.6550 1220.0000 265.6600 ;
      RECT 1214.5000 262.6550 1220.0000 265.6550 ;
      RECT 0.0000 262.6550 5.5000 265.6550 ;
      RECT 0.0000 260.6550 1220.0000 262.6550 ;
      RECT 1218.5000 257.6550 1220.0000 260.6550 ;
      RECT 0.0000 257.6550 1.5000 260.6550 ;
      RECT 0.0000 257.6500 1220.0000 257.6550 ;
      RECT 1214.5000 254.6500 1220.0000 257.6500 ;
      RECT 0.0000 254.6500 5.5000 257.6500 ;
      RECT 0.0000 252.6500 1220.0000 254.6500 ;
      RECT 1218.5000 249.6500 1220.0000 252.6500 ;
      RECT 0.0000 249.6500 1.5000 252.6500 ;
      RECT 0.0000 249.6450 1220.0000 249.6500 ;
      RECT 1214.5000 246.6450 1220.0000 249.6450 ;
      RECT 0.0000 246.6450 5.5000 249.6450 ;
      RECT 0.0000 244.6450 1220.0000 246.6450 ;
      RECT 1218.5000 241.6450 1220.0000 244.6450 ;
      RECT 0.0000 241.6450 1.5000 244.6450 ;
      RECT 0.0000 241.6400 1220.0000 241.6450 ;
      RECT 1214.5000 238.6400 1220.0000 241.6400 ;
      RECT 0.0000 238.6400 5.5000 241.6400 ;
      RECT 0.0000 236.6400 1220.0000 238.6400 ;
      RECT 1218.5000 233.6400 1220.0000 236.6400 ;
      RECT 0.0000 233.6400 1.5000 236.6400 ;
      RECT 0.0000 233.6350 1220.0000 233.6400 ;
      RECT 1214.5000 230.6350 1220.0000 233.6350 ;
      RECT 0.0000 230.6350 5.5000 233.6350 ;
      RECT 0.0000 228.6350 1220.0000 230.6350 ;
      RECT 1218.5000 225.6350 1220.0000 228.6350 ;
      RECT 0.0000 225.6350 1.5000 228.6350 ;
      RECT 0.0000 225.6300 1220.0000 225.6350 ;
      RECT 1214.5000 222.6300 1220.0000 225.6300 ;
      RECT 0.0000 222.6300 5.5000 225.6300 ;
      RECT 0.0000 220.6300 1220.0000 222.6300 ;
      RECT 1218.5000 217.6300 1220.0000 220.6300 ;
      RECT 0.0000 217.6300 1.5000 220.6300 ;
      RECT 0.0000 217.6250 1220.0000 217.6300 ;
      RECT 1214.5000 214.6250 1220.0000 217.6250 ;
      RECT 0.0000 214.6250 5.5000 217.6250 ;
      RECT 0.0000 212.6250 1220.0000 214.6250 ;
      RECT 1218.5000 209.6250 1220.0000 212.6250 ;
      RECT 0.0000 209.6250 1.5000 212.6250 ;
      RECT 0.0000 209.6200 1220.0000 209.6250 ;
      RECT 1214.5000 206.6200 1220.0000 209.6200 ;
      RECT 0.0000 206.6200 5.5000 209.6200 ;
      RECT 0.0000 204.6200 1220.0000 206.6200 ;
      RECT 1218.5000 201.6200 1220.0000 204.6200 ;
      RECT 0.0000 201.6200 1.5000 204.6200 ;
      RECT 0.0000 201.6150 1220.0000 201.6200 ;
      RECT 1214.5000 198.6150 1220.0000 201.6150 ;
      RECT 0.0000 198.6150 5.5000 201.6150 ;
      RECT 0.0000 196.6150 1220.0000 198.6150 ;
      RECT 1218.5000 193.6150 1220.0000 196.6150 ;
      RECT 0.0000 193.6150 1.5000 196.6150 ;
      RECT 0.0000 193.6100 1220.0000 193.6150 ;
      RECT 1214.5000 190.6100 1220.0000 193.6100 ;
      RECT 0.0000 190.6100 5.5000 193.6100 ;
      RECT 0.0000 188.6100 1220.0000 190.6100 ;
      RECT 1218.5000 185.6100 1220.0000 188.6100 ;
      RECT 0.0000 185.6100 1.5000 188.6100 ;
      RECT 0.0000 185.6050 1220.0000 185.6100 ;
      RECT 1214.5000 182.6050 1220.0000 185.6050 ;
      RECT 0.0000 182.6050 5.5000 185.6050 ;
      RECT 0.0000 180.6050 1220.0000 182.6050 ;
      RECT 1218.5000 177.6050 1220.0000 180.6050 ;
      RECT 0.0000 177.6050 1.5000 180.6050 ;
      RECT 0.0000 177.6000 1220.0000 177.6050 ;
      RECT 1214.5000 174.6000 1220.0000 177.6000 ;
      RECT 0.0000 174.6000 5.5000 177.6000 ;
      RECT 0.0000 172.6000 1220.0000 174.6000 ;
      RECT 1218.5000 169.6000 1220.0000 172.6000 ;
      RECT 0.0000 169.6000 1.5000 172.6000 ;
      RECT 0.0000 169.5950 1220.0000 169.6000 ;
      RECT 1214.5000 166.5950 1220.0000 169.5950 ;
      RECT 0.0000 166.5950 5.5000 169.5950 ;
      RECT 0.0000 164.5950 1220.0000 166.5950 ;
      RECT 1218.5000 161.5950 1220.0000 164.5950 ;
      RECT 0.0000 161.5950 1.5000 164.5950 ;
      RECT 0.0000 161.5900 1220.0000 161.5950 ;
      RECT 1214.5000 158.5900 1220.0000 161.5900 ;
      RECT 0.0000 158.5900 5.5000 161.5900 ;
      RECT 0.0000 156.5900 1220.0000 158.5900 ;
      RECT 1218.5000 153.5900 1220.0000 156.5900 ;
      RECT 0.0000 153.5900 1.5000 156.5900 ;
      RECT 0.0000 153.5850 1220.0000 153.5900 ;
      RECT 1214.5000 150.5850 1220.0000 153.5850 ;
      RECT 0.0000 150.5850 5.5000 153.5850 ;
      RECT 0.0000 148.5850 1220.0000 150.5850 ;
      RECT 1218.5000 145.5850 1220.0000 148.5850 ;
      RECT 0.0000 145.5850 1.5000 148.5850 ;
      RECT 0.0000 145.5800 1220.0000 145.5850 ;
      RECT 1214.5000 142.5800 1220.0000 145.5800 ;
      RECT 0.0000 142.5800 5.5000 145.5800 ;
      RECT 0.0000 140.5800 1220.0000 142.5800 ;
      RECT 1218.5000 137.5800 1220.0000 140.5800 ;
      RECT 0.0000 137.5800 1.5000 140.5800 ;
      RECT 0.0000 137.5750 1220.0000 137.5800 ;
      RECT 1214.5000 134.5750 1220.0000 137.5750 ;
      RECT 0.0000 134.5750 5.5000 137.5750 ;
      RECT 0.0000 132.5750 1220.0000 134.5750 ;
      RECT 1218.5000 129.5750 1220.0000 132.5750 ;
      RECT 0.0000 129.5750 1.5000 132.5750 ;
      RECT 0.0000 129.5700 1220.0000 129.5750 ;
      RECT 1214.5000 126.5700 1220.0000 129.5700 ;
      RECT 0.0000 126.5700 5.5000 129.5700 ;
      RECT 0.0000 124.5700 1220.0000 126.5700 ;
      RECT 1218.5000 121.5700 1220.0000 124.5700 ;
      RECT 0.0000 121.5700 1.5000 124.5700 ;
      RECT 0.0000 121.5650 1220.0000 121.5700 ;
      RECT 1214.5000 118.5650 1220.0000 121.5650 ;
      RECT 0.0000 118.5650 5.5000 121.5650 ;
      RECT 0.0000 116.5650 1220.0000 118.5650 ;
      RECT 1218.5000 113.5650 1220.0000 116.5650 ;
      RECT 0.0000 113.5650 1.5000 116.5650 ;
      RECT 0.0000 113.5600 1220.0000 113.5650 ;
      RECT 1214.5000 110.5600 1220.0000 113.5600 ;
      RECT 0.0000 110.5600 5.5000 113.5600 ;
      RECT 0.0000 108.5600 1220.0000 110.5600 ;
      RECT 1218.5000 105.5600 1220.0000 108.5600 ;
      RECT 0.0000 105.5600 1.5000 108.5600 ;
      RECT 0.0000 105.5550 1220.0000 105.5600 ;
      RECT 1214.5000 102.5550 1220.0000 105.5550 ;
      RECT 0.0000 102.5550 5.5000 105.5550 ;
      RECT 0.0000 100.5550 1220.0000 102.5550 ;
      RECT 1218.5000 97.5550 1220.0000 100.5550 ;
      RECT 0.0000 97.5550 1.5000 100.5550 ;
      RECT 0.0000 97.5500 1220.0000 97.5550 ;
      RECT 1214.5000 94.5500 1220.0000 97.5500 ;
      RECT 0.0000 94.5500 5.5000 97.5500 ;
      RECT 0.0000 92.5500 1220.0000 94.5500 ;
      RECT 1218.5000 89.5500 1220.0000 92.5500 ;
      RECT 0.0000 89.5500 1.5000 92.5500 ;
      RECT 0.0000 89.5450 1220.0000 89.5500 ;
      RECT 1214.5000 86.5450 1220.0000 89.5450 ;
      RECT 0.0000 86.5450 5.5000 89.5450 ;
      RECT 0.0000 84.5450 1220.0000 86.5450 ;
      RECT 1218.5000 81.5450 1220.0000 84.5450 ;
      RECT 0.0000 81.5450 1.5000 84.5450 ;
      RECT 0.0000 81.5400 1220.0000 81.5450 ;
      RECT 1214.5000 78.5400 1220.0000 81.5400 ;
      RECT 0.0000 78.5400 5.5000 81.5400 ;
      RECT 0.0000 76.5400 1220.0000 78.5400 ;
      RECT 1218.5000 73.5400 1220.0000 76.5400 ;
      RECT 0.0000 73.5400 1.5000 76.5400 ;
      RECT 0.0000 73.5350 1220.0000 73.5400 ;
      RECT 1214.5000 70.5350 1220.0000 73.5350 ;
      RECT 0.0000 70.5350 5.5000 73.5350 ;
      RECT 0.0000 68.5350 1220.0000 70.5350 ;
      RECT 1218.5000 65.5350 1220.0000 68.5350 ;
      RECT 0.0000 65.5350 1.5000 68.5350 ;
      RECT 0.0000 65.5300 1220.0000 65.5350 ;
      RECT 1214.5000 62.5300 1220.0000 65.5300 ;
      RECT 0.0000 62.5300 5.5000 65.5300 ;
      RECT 0.0000 60.5300 1220.0000 62.5300 ;
      RECT 1218.5000 57.5300 1220.0000 60.5300 ;
      RECT 0.0000 57.5300 1.5000 60.5300 ;
      RECT 0.0000 57.5250 1220.0000 57.5300 ;
      RECT 1214.5000 54.5250 1220.0000 57.5250 ;
      RECT 0.0000 54.5250 5.5000 57.5250 ;
      RECT 0.0000 52.5250 1220.0000 54.5250 ;
      RECT 1218.5000 49.5250 1220.0000 52.5250 ;
      RECT 0.0000 49.5250 1.5000 52.5250 ;
      RECT 0.0000 49.5200 1220.0000 49.5250 ;
      RECT 1214.5000 46.5200 1220.0000 49.5200 ;
      RECT 0.0000 46.5200 5.5000 49.5200 ;
      RECT 0.0000 44.5200 1220.0000 46.5200 ;
      RECT 1218.5000 41.5200 1220.0000 44.5200 ;
      RECT 0.0000 41.5200 1.5000 44.5200 ;
      RECT 0.0000 41.5150 1220.0000 41.5200 ;
      RECT 1214.5000 38.5150 1220.0000 41.5150 ;
      RECT 0.0000 38.5150 5.5000 41.5150 ;
      RECT 0.0000 36.5150 1220.0000 38.5150 ;
      RECT 1218.5000 33.5150 1220.0000 36.5150 ;
      RECT 0.0000 33.5150 1.5000 36.5150 ;
      RECT 0.0000 33.5100 1220.0000 33.5150 ;
      RECT 1214.5000 30.5100 1220.0000 33.5100 ;
      RECT 0.0000 30.5100 5.5000 33.5100 ;
      RECT 0.0000 28.5100 1220.0000 30.5100 ;
      RECT 1218.5000 25.5100 1220.0000 28.5100 ;
      RECT 0.0000 25.5100 1.5000 28.5100 ;
      RECT 0.0000 25.5050 1220.0000 25.5100 ;
      RECT 1214.5000 22.5050 1220.0000 25.5050 ;
      RECT 0.0000 22.5050 5.5000 25.5050 ;
      RECT 0.0000 20.5050 1220.0000 22.5050 ;
      RECT 1218.5000 17.5050 1220.0000 20.5050 ;
      RECT 0.0000 17.5050 1.5000 20.5050 ;
      RECT 0.0000 17.5000 1220.0000 17.5050 ;
      RECT 1214.5000 14.5000 1220.0000 17.5000 ;
      RECT 0.0000 14.5000 5.5000 17.5000 ;
      RECT 0.0000 12.5000 1220.0000 14.5000 ;
      RECT 1218.5000 9.5000 1220.0000 12.5000 ;
      RECT 0.0000 9.5000 1.5000 12.5000 ;
      RECT 0.0000 0.0000 1220.0000 9.5000 ;
  END
END core

END LIBRARY
