##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Tue Mar 18 21:26:34 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16_160b
  CLASS BLOCK ;
  SIZE 670.0000 BY 670.0000 ;
  FOREIGN sram_w16_160b 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 342.7500 0.5200 342.8500 ;
    END
  END CLK
  PIN D[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 652.8500 0.0000 652.9500 0.5200 ;
    END
  END D[159]
  PIN D[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 648.8500 0.0000 648.9500 0.5200 ;
    END
  END D[158]
  PIN D[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 644.8500 0.0000 644.9500 0.5200 ;
    END
  END D[157]
  PIN D[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 640.8500 0.0000 640.9500 0.5200 ;
    END
  END D[156]
  PIN D[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 636.8500 0.0000 636.9500 0.5200 ;
    END
  END D[155]
  PIN D[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 632.8500 0.0000 632.9500 0.5200 ;
    END
  END D[154]
  PIN D[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 628.8500 0.0000 628.9500 0.5200 ;
    END
  END D[153]
  PIN D[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 624.8500 0.0000 624.9500 0.5200 ;
    END
  END D[152]
  PIN D[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 620.8500 0.0000 620.9500 0.5200 ;
    END
  END D[151]
  PIN D[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 616.8500 0.0000 616.9500 0.5200 ;
    END
  END D[150]
  PIN D[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 612.8500 0.0000 612.9500 0.5200 ;
    END
  END D[149]
  PIN D[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 608.8500 0.0000 608.9500 0.5200 ;
    END
  END D[148]
  PIN D[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 604.8500 0.0000 604.9500 0.5200 ;
    END
  END D[147]
  PIN D[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 600.8500 0.0000 600.9500 0.5200 ;
    END
  END D[146]
  PIN D[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 596.8500 0.0000 596.9500 0.5200 ;
    END
  END D[145]
  PIN D[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 592.8500 0.0000 592.9500 0.5200 ;
    END
  END D[144]
  PIN D[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 588.8500 0.0000 588.9500 0.5200 ;
    END
  END D[143]
  PIN D[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 584.8500 0.0000 584.9500 0.5200 ;
    END
  END D[142]
  PIN D[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 580.8500 0.0000 580.9500 0.5200 ;
    END
  END D[141]
  PIN D[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 576.8500 0.0000 576.9500 0.5200 ;
    END
  END D[140]
  PIN D[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 572.8500 0.0000 572.9500 0.5200 ;
    END
  END D[139]
  PIN D[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 568.8500 0.0000 568.9500 0.5200 ;
    END
  END D[138]
  PIN D[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 564.8500 0.0000 564.9500 0.5200 ;
    END
  END D[137]
  PIN D[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 560.8500 0.0000 560.9500 0.5200 ;
    END
  END D[136]
  PIN D[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 556.8500 0.0000 556.9500 0.5200 ;
    END
  END D[135]
  PIN D[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 552.8500 0.0000 552.9500 0.5200 ;
    END
  END D[134]
  PIN D[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 548.8500 0.0000 548.9500 0.5200 ;
    END
  END D[133]
  PIN D[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 544.8500 0.0000 544.9500 0.5200 ;
    END
  END D[132]
  PIN D[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 540.8500 0.0000 540.9500 0.5200 ;
    END
  END D[131]
  PIN D[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.8500 0.0000 536.9500 0.5200 ;
    END
  END D[130]
  PIN D[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 532.8500 0.0000 532.9500 0.5200 ;
    END
  END D[129]
  PIN D[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 528.8500 0.0000 528.9500 0.5200 ;
    END
  END D[128]
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 524.8500 0.0000 524.9500 0.5200 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 520.8500 0.0000 520.9500 0.5200 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 516.8500 0.0000 516.9500 0.5200 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 512.8500 0.0000 512.9500 0.5200 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 508.8500 0.0000 508.9500 0.5200 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 504.8500 0.0000 504.9500 0.5200 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 500.8500 0.0000 500.9500 0.5200 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 496.8500 0.0000 496.9500 0.5200 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 492.8500 0.0000 492.9500 0.5200 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 488.8500 0.0000 488.9500 0.5200 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 484.8500 0.0000 484.9500 0.5200 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 480.8500 0.0000 480.9500 0.5200 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 476.8500 0.0000 476.9500 0.5200 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 472.8500 0.0000 472.9500 0.5200 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 468.8500 0.0000 468.9500 0.5200 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 464.8500 0.0000 464.9500 0.5200 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 460.8500 0.0000 460.9500 0.5200 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.8500 0.0000 456.9500 0.5200 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.8500 0.0000 452.9500 0.5200 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.8500 0.0000 448.9500 0.5200 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.8500 0.0000 444.9500 0.5200 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.8500 0.0000 440.9500 0.5200 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.8500 0.0000 436.9500 0.5200 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.8500 0.0000 432.9500 0.5200 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.8500 0.0000 428.9500 0.5200 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.8500 0.0000 424.9500 0.5200 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.8500 0.0000 420.9500 0.5200 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 416.8500 0.0000 416.9500 0.5200 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.8500 0.0000 412.9500 0.5200 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.8500 0.0000 408.9500 0.5200 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.8500 0.0000 404.9500 0.5200 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.8500 0.0000 400.9500 0.5200 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.8500 0.0000 396.9500 0.5200 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.8500 0.0000 392.9500 0.5200 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.8500 0.0000 388.9500 0.5200 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.8500 0.0000 384.9500 0.5200 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.8500 0.0000 380.9500 0.5200 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.8500 0.0000 376.9500 0.5200 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.8500 0.0000 372.9500 0.5200 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.8500 0.0000 368.9500 0.5200 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.8500 0.0000 364.9500 0.5200 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.8500 0.0000 360.9500 0.5200 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.8500 0.0000 356.9500 0.5200 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.8500 0.0000 352.9500 0.5200 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.8500 0.0000 348.9500 0.5200 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.8500 0.0000 344.9500 0.5200 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.8500 0.0000 340.9500 0.5200 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.8500 0.0000 336.9500 0.5200 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.8500 0.0000 332.9500 0.5200 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.8500 0.0000 328.9500 0.5200 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.8500 0.0000 324.9500 0.5200 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.8500 0.0000 320.9500 0.5200 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.8500 0.0000 316.9500 0.5200 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.8500 0.0000 312.9500 0.5200 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.8500 0.0000 308.9500 0.5200 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 304.8500 0.0000 304.9500 0.5200 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.8500 0.0000 300.9500 0.5200 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 296.8500 0.0000 296.9500 0.5200 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 292.8500 0.0000 292.9500 0.5200 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.8500 0.0000 288.9500 0.5200 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284.8500 0.0000 284.9500 0.5200 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.8500 0.0000 280.9500 0.5200 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 276.8500 0.0000 276.9500 0.5200 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 272.8500 0.0000 272.9500 0.5200 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.8500 0.0000 268.9500 0.5200 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 264.8500 0.0000 264.9500 0.5200 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.8500 0.0000 260.9500 0.5200 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.8500 0.0000 256.9500 0.5200 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.8500 0.0000 252.9500 0.5200 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.8500 0.0000 248.9500 0.5200 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.8500 0.0000 244.9500 0.5200 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.8500 0.0000 240.9500 0.5200 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 236.8500 0.0000 236.9500 0.5200 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.8500 0.0000 232.9500 0.5200 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.8500 0.0000 228.9500 0.5200 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.8500 0.0000 224.9500 0.5200 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.8500 0.0000 220.9500 0.5200 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.8500 0.0000 216.9500 0.5200 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.8500 0.0000 212.9500 0.5200 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.8500 0.0000 208.9500 0.5200 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.8500 0.0000 204.9500 0.5200 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.8500 0.0000 200.9500 0.5200 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.8500 0.0000 196.9500 0.5200 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.8500 0.0000 192.9500 0.5200 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.8500 0.0000 188.9500 0.5200 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.8500 0.0000 184.9500 0.5200 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.8500 0.0000 180.9500 0.5200 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.8500 0.0000 176.9500 0.5200 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.8500 0.0000 172.9500 0.5200 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.8500 0.0000 168.9500 0.5200 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.8500 0.0000 164.9500 0.5200 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.8500 0.0000 160.9500 0.5200 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.8500 0.0000 156.9500 0.5200 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.8500 0.0000 152.9500 0.5200 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.8500 0.0000 148.9500 0.5200 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.8500 0.0000 144.9500 0.5200 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.8500 0.0000 140.9500 0.5200 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.8500 0.0000 136.9500 0.5200 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.8500 0.0000 132.9500 0.5200 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.8500 0.0000 128.9500 0.5200 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.8500 0.0000 124.9500 0.5200 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.8500 0.0000 120.9500 0.5200 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.8500 0.0000 116.9500 0.5200 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.8500 0.0000 112.9500 0.5200 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.8500 0.0000 108.9500 0.5200 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.8500 0.0000 104.9500 0.5200 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.8500 0.0000 100.9500 0.5200 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.8500 0.0000 96.9500 0.5200 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.8500 0.0000 92.9500 0.5200 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.8500 0.0000 88.9500 0.5200 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.8500 0.0000 84.9500 0.5200 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.8500 0.0000 80.9500 0.5200 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.8500 0.0000 76.9500 0.5200 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.8500 0.0000 72.9500 0.5200 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.8500 0.0000 68.9500 0.5200 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.8500 0.0000 64.9500 0.5200 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.8500 0.0000 60.9500 0.5200 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.8500 0.0000 56.9500 0.5200 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.8500 0.0000 52.9500 0.5200 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.8500 0.0000 48.9500 0.5200 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.8500 0.0000 44.9500 0.5200 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.8500 0.0000 40.9500 0.5200 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.8500 0.0000 36.9500 0.5200 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.8500 0.0000 32.9500 0.5200 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.8500 0.0000 28.9500 0.5200 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.8500 0.0000 24.9500 0.5200 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.8500 0.0000 20.9500 0.5200 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.8500 0.0000 16.9500 0.5200 ;
    END
  END D[0]
  PIN Q[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 652.8500 669.4800 652.9500 670.0000 ;
    END
  END Q[159]
  PIN Q[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 648.8500 669.4800 648.9500 670.0000 ;
    END
  END Q[158]
  PIN Q[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 644.8500 669.4800 644.9500 670.0000 ;
    END
  END Q[157]
  PIN Q[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 640.8500 669.4800 640.9500 670.0000 ;
    END
  END Q[156]
  PIN Q[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 636.8500 669.4800 636.9500 670.0000 ;
    END
  END Q[155]
  PIN Q[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 632.8500 669.4800 632.9500 670.0000 ;
    END
  END Q[154]
  PIN Q[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 628.8500 669.4800 628.9500 670.0000 ;
    END
  END Q[153]
  PIN Q[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 624.8500 669.4800 624.9500 670.0000 ;
    END
  END Q[152]
  PIN Q[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 620.8500 669.4800 620.9500 670.0000 ;
    END
  END Q[151]
  PIN Q[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 616.8500 669.4800 616.9500 670.0000 ;
    END
  END Q[150]
  PIN Q[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 612.8500 669.4800 612.9500 670.0000 ;
    END
  END Q[149]
  PIN Q[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 608.8500 669.4800 608.9500 670.0000 ;
    END
  END Q[148]
  PIN Q[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 604.8500 669.4800 604.9500 670.0000 ;
    END
  END Q[147]
  PIN Q[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 600.8500 669.4800 600.9500 670.0000 ;
    END
  END Q[146]
  PIN Q[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 596.8500 669.4800 596.9500 670.0000 ;
    END
  END Q[145]
  PIN Q[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 592.8500 669.4800 592.9500 670.0000 ;
    END
  END Q[144]
  PIN Q[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 588.8500 669.4800 588.9500 670.0000 ;
    END
  END Q[143]
  PIN Q[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 584.8500 669.4800 584.9500 670.0000 ;
    END
  END Q[142]
  PIN Q[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 580.8500 669.4800 580.9500 670.0000 ;
    END
  END Q[141]
  PIN Q[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 576.8500 669.4800 576.9500 670.0000 ;
    END
  END Q[140]
  PIN Q[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 572.8500 669.4800 572.9500 670.0000 ;
    END
  END Q[139]
  PIN Q[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 568.8500 669.4800 568.9500 670.0000 ;
    END
  END Q[138]
  PIN Q[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 564.8500 669.4800 564.9500 670.0000 ;
    END
  END Q[137]
  PIN Q[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 560.8500 669.4800 560.9500 670.0000 ;
    END
  END Q[136]
  PIN Q[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 556.8500 669.4800 556.9500 670.0000 ;
    END
  END Q[135]
  PIN Q[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 552.8500 669.4800 552.9500 670.0000 ;
    END
  END Q[134]
  PIN Q[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 548.8500 669.4800 548.9500 670.0000 ;
    END
  END Q[133]
  PIN Q[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 544.8500 669.4800 544.9500 670.0000 ;
    END
  END Q[132]
  PIN Q[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 540.8500 669.4800 540.9500 670.0000 ;
    END
  END Q[131]
  PIN Q[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.8500 669.4800 536.9500 670.0000 ;
    END
  END Q[130]
  PIN Q[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 532.8500 669.4800 532.9500 670.0000 ;
    END
  END Q[129]
  PIN Q[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 528.8500 669.4800 528.9500 670.0000 ;
    END
  END Q[128]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 524.8500 669.4800 524.9500 670.0000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 520.8500 669.4800 520.9500 670.0000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 516.8500 669.4800 516.9500 670.0000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 512.8500 669.4800 512.9500 670.0000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 508.8500 669.4800 508.9500 670.0000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 504.8500 669.4800 504.9500 670.0000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 500.8500 669.4800 500.9500 670.0000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 496.8500 669.4800 496.9500 670.0000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 492.8500 669.4800 492.9500 670.0000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 488.8500 669.4800 488.9500 670.0000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 484.8500 669.4800 484.9500 670.0000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 480.8500 669.4800 480.9500 670.0000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 476.8500 669.4800 476.9500 670.0000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 472.8500 669.4800 472.9500 670.0000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 468.8500 669.4800 468.9500 670.0000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 464.8500 669.4800 464.9500 670.0000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 460.8500 669.4800 460.9500 670.0000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.8500 669.4800 456.9500 670.0000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.8500 669.4800 452.9500 670.0000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.8500 669.4800 448.9500 670.0000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.8500 669.4800 444.9500 670.0000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.8500 669.4800 440.9500 670.0000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.8500 669.4800 436.9500 670.0000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.8500 669.4800 432.9500 670.0000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.8500 669.4800 428.9500 670.0000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.8500 669.4800 424.9500 670.0000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.8500 669.4800 420.9500 670.0000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 416.8500 669.4800 416.9500 670.0000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.8500 669.4800 412.9500 670.0000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.8500 669.4800 408.9500 670.0000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.8500 669.4800 404.9500 670.0000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.8500 669.4800 400.9500 670.0000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.8500 669.4800 396.9500 670.0000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.8500 669.4800 392.9500 670.0000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.8500 669.4800 388.9500 670.0000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.8500 669.4800 384.9500 670.0000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.8500 669.4800 380.9500 670.0000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.8500 669.4800 376.9500 670.0000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.8500 669.4800 372.9500 670.0000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.8500 669.4800 368.9500 670.0000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.8500 669.4800 364.9500 670.0000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.8500 669.4800 360.9500 670.0000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.8500 669.4800 356.9500 670.0000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.8500 669.4800 352.9500 670.0000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.8500 669.4800 348.9500 670.0000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.8500 669.4800 344.9500 670.0000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.8500 669.4800 340.9500 670.0000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.8500 669.4800 336.9500 670.0000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.8500 669.4800 332.9500 670.0000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.8500 669.4800 328.9500 670.0000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.8500 669.4800 324.9500 670.0000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.8500 669.4800 320.9500 670.0000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.8500 669.4800 316.9500 670.0000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.8500 669.4800 312.9500 670.0000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.8500 669.4800 308.9500 670.0000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 304.8500 669.4800 304.9500 670.0000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.8500 669.4800 300.9500 670.0000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 296.8500 669.4800 296.9500 670.0000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 292.8500 669.4800 292.9500 670.0000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.8500 669.4800 288.9500 670.0000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284.8500 669.4800 284.9500 670.0000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.8500 669.4800 280.9500 670.0000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 276.8500 669.4800 276.9500 670.0000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 272.8500 669.4800 272.9500 670.0000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.8500 669.4800 268.9500 670.0000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 264.8500 669.4800 264.9500 670.0000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.8500 669.4800 260.9500 670.0000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.8500 669.4800 256.9500 670.0000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.8500 669.4800 252.9500 670.0000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.8500 669.4800 248.9500 670.0000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.8500 669.4800 244.9500 670.0000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.8500 669.4800 240.9500 670.0000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 236.8500 669.4800 236.9500 670.0000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.8500 669.4800 232.9500 670.0000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.8500 669.4800 228.9500 670.0000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.8500 669.4800 224.9500 670.0000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.8500 669.4800 220.9500 670.0000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.8500 669.4800 216.9500 670.0000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.8500 669.4800 212.9500 670.0000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.8500 669.4800 208.9500 670.0000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.8500 669.4800 204.9500 670.0000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.8500 669.4800 200.9500 670.0000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.8500 669.4800 196.9500 670.0000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.8500 669.4800 192.9500 670.0000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.8500 669.4800 188.9500 670.0000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.8500 669.4800 184.9500 670.0000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.8500 669.4800 180.9500 670.0000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.8500 669.4800 176.9500 670.0000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.8500 669.4800 172.9500 670.0000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.8500 669.4800 168.9500 670.0000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.8500 669.4800 164.9500 670.0000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.8500 669.4800 160.9500 670.0000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.8500 669.4800 156.9500 670.0000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.8500 669.4800 152.9500 670.0000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.8500 669.4800 148.9500 670.0000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.8500 669.4800 144.9500 670.0000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.8500 669.4800 140.9500 670.0000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.8500 669.4800 136.9500 670.0000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.8500 669.4800 132.9500 670.0000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.8500 669.4800 128.9500 670.0000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.8500 669.4800 124.9500 670.0000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.8500 669.4800 120.9500 670.0000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.8500 669.4800 116.9500 670.0000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.8500 669.4800 112.9500 670.0000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.8500 669.4800 108.9500 670.0000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.8500 669.4800 104.9500 670.0000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.8500 669.4800 100.9500 670.0000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.8500 669.4800 96.9500 670.0000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.8500 669.4800 92.9500 670.0000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.8500 669.4800 88.9500 670.0000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.8500 669.4800 84.9500 670.0000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.8500 669.4800 80.9500 670.0000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.8500 669.4800 76.9500 670.0000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.8500 669.4800 72.9500 670.0000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.8500 669.4800 68.9500 670.0000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.8500 669.4800 64.9500 670.0000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.8500 669.4800 60.9500 670.0000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.8500 669.4800 56.9500 670.0000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.8500 669.4800 52.9500 670.0000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.8500 669.4800 48.9500 670.0000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.8500 669.4800 44.9500 670.0000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.8500 669.4800 40.9500 670.0000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.8500 669.4800 36.9500 670.0000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.8500 669.4800 32.9500 670.0000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.8500 669.4800 28.9500 670.0000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.8500 669.4800 24.9500 670.0000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.8500 669.4800 20.9500 670.0000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.8500 669.4800 16.9500 670.0000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 338.7500 0.5200 338.8500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 346.7500 0.5200 346.8500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 334.7500 0.5200 334.8500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 330.7500 0.5200 330.8500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 326.7500 0.5200 326.8500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 322.7500 0.5200 322.8500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 83.3500 10.0000 85.3500 660.0000 ;
        RECT 75.2000 10.0000 77.2000 660.0000 ;
        RECT 67.0500 10.0000 69.0500 660.0000 ;
        RECT 58.9000 10.0000 60.9000 660.0000 ;
        RECT 50.7500 10.0000 52.7500 660.0000 ;
        RECT 42.6000 10.0000 44.6000 660.0000 ;
        RECT 34.4500 10.0000 36.4500 660.0000 ;
        RECT 26.3000 10.0000 28.3000 660.0000 ;
        RECT 18.1500 10.0000 20.1500 660.0000 ;
        RECT 10.0000 10.0000 12.0000 660.0000 ;
        RECT 164.8500 10.0000 166.8500 660.0000 ;
        RECT 156.7000 10.0000 158.7000 660.0000 ;
        RECT 148.5500 10.0000 150.5500 660.0000 ;
        RECT 140.4000 10.0000 142.4000 660.0000 ;
        RECT 132.2500 10.0000 134.2500 660.0000 ;
        RECT 124.1000 10.0000 126.1000 660.0000 ;
        RECT 115.9500 10.0000 117.9500 660.0000 ;
        RECT 107.8000 10.0000 109.8000 660.0000 ;
        RECT 99.6500 10.0000 101.6500 660.0000 ;
        RECT 91.5000 10.0000 93.5000 660.0000 ;
        RECT 246.3500 10.0000 248.3500 660.0000 ;
        RECT 238.2000 10.0000 240.2000 660.0000 ;
        RECT 230.0500 10.0000 232.0500 660.0000 ;
        RECT 221.9000 10.0000 223.9000 660.0000 ;
        RECT 213.7500 10.0000 215.7500 660.0000 ;
        RECT 205.6000 10.0000 207.6000 660.0000 ;
        RECT 197.4500 10.0000 199.4500 660.0000 ;
        RECT 189.3000 10.0000 191.3000 660.0000 ;
        RECT 181.1500 10.0000 183.1500 660.0000 ;
        RECT 173.0000 10.0000 175.0000 660.0000 ;
        RECT 327.8500 10.0000 329.8500 660.0000 ;
        RECT 319.7000 10.0000 321.7000 660.0000 ;
        RECT 311.5500 10.0000 313.5500 660.0000 ;
        RECT 303.4000 10.0000 305.4000 660.0000 ;
        RECT 295.2500 10.0000 297.2500 660.0000 ;
        RECT 287.1000 10.0000 289.1000 660.0000 ;
        RECT 278.9500 10.0000 280.9500 660.0000 ;
        RECT 270.8000 10.0000 272.8000 660.0000 ;
        RECT 254.5000 10.0000 256.5000 660.0000 ;
        RECT 262.6500 10.0000 264.6500 660.0000 ;
        RECT 417.5000 10.0000 419.5000 660.0000 ;
        RECT 336.0000 10.0000 338.0000 660.0000 ;
        RECT 344.1500 10.0000 346.1500 660.0000 ;
        RECT 352.3000 10.0000 354.3000 660.0000 ;
        RECT 360.4500 10.0000 362.4500 660.0000 ;
        RECT 368.6000 10.0000 370.6000 660.0000 ;
        RECT 376.7500 10.0000 378.7500 660.0000 ;
        RECT 384.9000 10.0000 386.9000 660.0000 ;
        RECT 393.0500 10.0000 395.0500 660.0000 ;
        RECT 401.2000 10.0000 403.2000 660.0000 ;
        RECT 409.3500 10.0000 411.3500 660.0000 ;
        RECT 425.6500 10.0000 427.6500 660.0000 ;
        RECT 433.8000 10.0000 435.8000 660.0000 ;
        RECT 441.9500 10.0000 443.9500 660.0000 ;
        RECT 450.1000 10.0000 452.1000 660.0000 ;
        RECT 458.2500 10.0000 460.2500 660.0000 ;
        RECT 466.4000 10.0000 468.4000 660.0000 ;
        RECT 474.5500 10.0000 476.5500 660.0000 ;
        RECT 482.7000 10.0000 484.7000 660.0000 ;
        RECT 490.8500 10.0000 492.8500 660.0000 ;
        RECT 499.0000 10.0000 501.0000 660.0000 ;
        RECT 580.5000 10.0000 582.5000 660.0000 ;
        RECT 507.1500 10.0000 509.1500 660.0000 ;
        RECT 515.3000 10.0000 517.3000 660.0000 ;
        RECT 523.4500 10.0000 525.4500 660.0000 ;
        RECT 531.6000 10.0000 533.6000 660.0000 ;
        RECT 539.7500 10.0000 541.7500 660.0000 ;
        RECT 547.9000 10.0000 549.9000 660.0000 ;
        RECT 556.0500 10.0000 558.0500 660.0000 ;
        RECT 564.2000 10.0000 566.2000 660.0000 ;
        RECT 572.3500 10.0000 574.3500 660.0000 ;
        RECT 653.8500 10.0000 655.8500 660.0000 ;
        RECT 645.7000 10.0000 647.7000 660.0000 ;
        RECT 637.5500 10.0000 639.5500 660.0000 ;
        RECT 629.4000 10.0000 631.4000 660.0000 ;
        RECT 621.2500 10.0000 623.2500 660.0000 ;
        RECT 613.1000 10.0000 615.1000 660.0000 ;
        RECT 604.9500 10.0000 606.9500 660.0000 ;
        RECT 596.8000 10.0000 598.8000 660.0000 ;
        RECT 588.6500 10.0000 590.6500 660.0000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 79.2000 10.0000 81.2000 660.0000 ;
        RECT 71.0500 10.0000 73.0500 660.0000 ;
        RECT 62.9000 10.0000 64.9000 660.0000 ;
        RECT 54.7500 10.0000 56.7500 660.0000 ;
        RECT 46.6000 10.0000 48.6000 660.0000 ;
        RECT 38.4500 10.0000 40.4500 660.0000 ;
        RECT 30.3000 10.0000 32.3000 660.0000 ;
        RECT 22.1500 10.0000 24.1500 660.0000 ;
        RECT 14.0000 10.0000 16.0000 660.0000 ;
        RECT 87.3500 10.0000 89.3500 660.0000 ;
        RECT 95.5000 10.0000 97.5000 660.0000 ;
        RECT 103.6500 10.0000 105.6500 660.0000 ;
        RECT 111.8000 10.0000 113.8000 660.0000 ;
        RECT 119.9500 10.0000 121.9500 660.0000 ;
        RECT 128.1000 10.0000 130.1000 660.0000 ;
        RECT 136.2500 10.0000 138.2500 660.0000 ;
        RECT 144.4000 10.0000 146.4000 660.0000 ;
        RECT 152.5500 10.0000 154.5500 660.0000 ;
        RECT 160.7000 10.0000 162.7000 660.0000 ;
        RECT 250.3500 10.0000 252.3500 660.0000 ;
        RECT 242.2000 10.0000 244.2000 660.0000 ;
        RECT 234.0500 10.0000 236.0500 660.0000 ;
        RECT 225.9000 10.0000 227.9000 660.0000 ;
        RECT 217.7500 10.0000 219.7500 660.0000 ;
        RECT 209.6000 10.0000 211.6000 660.0000 ;
        RECT 201.4500 10.0000 203.4500 660.0000 ;
        RECT 193.3000 10.0000 195.3000 660.0000 ;
        RECT 185.1500 10.0000 187.1500 660.0000 ;
        RECT 177.0000 10.0000 179.0000 660.0000 ;
        RECT 168.8500 10.0000 170.8500 660.0000 ;
        RECT 258.5000 10.0000 260.5000 660.0000 ;
        RECT 266.6500 10.0000 268.6500 660.0000 ;
        RECT 274.8000 10.0000 276.8000 660.0000 ;
        RECT 282.9500 10.0000 284.9500 660.0000 ;
        RECT 291.1000 10.0000 293.1000 660.0000 ;
        RECT 299.2500 10.0000 301.2500 660.0000 ;
        RECT 307.4000 10.0000 309.4000 660.0000 ;
        RECT 315.5500 10.0000 317.5500 660.0000 ;
        RECT 323.7000 10.0000 325.7000 660.0000 ;
        RECT 331.8500 10.0000 333.8500 660.0000 ;
        RECT 405.2000 10.0000 407.2000 660.0000 ;
        RECT 397.0500 10.0000 399.0500 660.0000 ;
        RECT 388.9000 10.0000 390.9000 660.0000 ;
        RECT 380.7500 10.0000 382.7500 660.0000 ;
        RECT 372.6000 10.0000 374.6000 660.0000 ;
        RECT 364.4500 10.0000 366.4500 660.0000 ;
        RECT 356.3000 10.0000 358.3000 660.0000 ;
        RECT 348.1500 10.0000 350.1500 660.0000 ;
        RECT 340.0000 10.0000 342.0000 660.0000 ;
        RECT 413.3500 10.0000 415.3500 660.0000 ;
        RECT 421.5000 10.0000 423.5000 660.0000 ;
        RECT 429.6500 10.0000 431.6500 660.0000 ;
        RECT 437.8000 10.0000 439.8000 660.0000 ;
        RECT 445.9500 10.0000 447.9500 660.0000 ;
        RECT 454.1000 10.0000 456.1000 660.0000 ;
        RECT 462.2500 10.0000 464.2500 660.0000 ;
        RECT 470.4000 10.0000 472.4000 660.0000 ;
        RECT 478.5500 10.0000 480.5500 660.0000 ;
        RECT 486.7000 10.0000 488.7000 660.0000 ;
        RECT 494.8500 10.0000 496.8500 660.0000 ;
        RECT 584.5000 10.0000 586.5000 660.0000 ;
        RECT 576.3500 10.0000 578.3500 660.0000 ;
        RECT 568.2000 10.0000 570.2000 660.0000 ;
        RECT 560.0500 10.0000 562.0500 660.0000 ;
        RECT 551.9000 10.0000 553.9000 660.0000 ;
        RECT 543.7500 10.0000 545.7500 660.0000 ;
        RECT 535.6000 10.0000 537.6000 660.0000 ;
        RECT 527.4500 10.0000 529.4500 660.0000 ;
        RECT 519.3000 10.0000 521.3000 660.0000 ;
        RECT 511.1500 10.0000 513.1500 660.0000 ;
        RECT 503.0000 10.0000 505.0000 660.0000 ;
        RECT 592.6500 10.0000 594.6500 660.0000 ;
        RECT 600.8000 10.0000 602.8000 660.0000 ;
        RECT 608.9500 10.0000 610.9500 660.0000 ;
        RECT 617.1000 10.0000 619.1000 660.0000 ;
        RECT 625.2500 10.0000 627.2500 660.0000 ;
        RECT 633.4000 10.0000 635.4000 660.0000 ;
        RECT 641.5500 10.0000 643.5500 660.0000 ;
        RECT 649.7000 10.0000 651.7000 660.0000 ;
        RECT 657.8500 10.0000 659.8500 660.0000 ;
        RECT 14.0000 9.8350 16.0000 10.1650 ;
        RECT 38.4500 9.8350 40.4500 10.1650 ;
        RECT 30.3000 9.8350 32.3000 10.1650 ;
        RECT 22.1500 9.8350 24.1500 10.1650 ;
        RECT 54.7500 9.8350 56.7500 10.1650 ;
        RECT 46.6000 9.8350 48.6000 10.1650 ;
        RECT 79.2000 9.8350 81.2000 10.1650 ;
        RECT 71.0500 9.8350 73.0500 10.1650 ;
        RECT 62.9000 9.8350 64.9000 10.1650 ;
        RECT 103.6500 9.8350 105.6500 10.1650 ;
        RECT 95.5000 9.8350 97.5000 10.1650 ;
        RECT 87.3500 9.8350 89.3500 10.1650 ;
        RECT 119.9500 9.8350 121.9500 10.1650 ;
        RECT 111.8000 9.8350 113.8000 10.1650 ;
        RECT 144.4000 9.8350 146.4000 10.1650 ;
        RECT 136.2500 9.8350 138.2500 10.1650 ;
        RECT 128.1000 9.8350 130.1000 10.1650 ;
        RECT 160.7000 9.8350 162.7000 10.1650 ;
        RECT 152.5500 9.8350 154.5500 10.1650 ;
        RECT 250.3500 9.8350 252.3500 10.1650 ;
        RECT 185.1500 9.8350 187.1500 10.1650 ;
        RECT 177.0000 9.8350 179.0000 10.1650 ;
        RECT 168.8500 9.8350 170.8500 10.1650 ;
        RECT 201.4500 9.8350 203.4500 10.1650 ;
        RECT 193.3000 9.8350 195.3000 10.1650 ;
        RECT 225.9000 9.8350 227.9000 10.1650 ;
        RECT 217.7500 9.8350 219.7500 10.1650 ;
        RECT 209.6000 9.8350 211.6000 10.1650 ;
        RECT 242.2000 9.8350 244.2000 10.1650 ;
        RECT 234.0500 9.8350 236.0500 10.1650 ;
        RECT 266.6500 9.8350 268.6500 10.1650 ;
        RECT 258.5000 9.8350 260.5000 10.1650 ;
        RECT 291.1000 9.8350 293.1000 10.1650 ;
        RECT 282.9500 9.8350 284.9500 10.1650 ;
        RECT 274.8000 9.8350 276.8000 10.1650 ;
        RECT 307.4000 9.8350 309.4000 10.1650 ;
        RECT 299.2500 9.8350 301.2500 10.1650 ;
        RECT 331.8500 9.8350 333.8500 10.1650 ;
        RECT 323.7000 9.8350 325.7000 10.1650 ;
        RECT 315.5500 9.8350 317.5500 10.1650 ;
        RECT 348.1500 9.8350 350.1500 10.1650 ;
        RECT 340.0000 9.8350 342.0000 10.1650 ;
        RECT 372.6000 9.8350 374.6000 10.1650 ;
        RECT 364.4500 9.8350 366.4500 10.1650 ;
        RECT 356.3000 9.8350 358.3000 10.1650 ;
        RECT 397.0500 9.8350 399.0500 10.1650 ;
        RECT 388.9000 9.8350 390.9000 10.1650 ;
        RECT 380.7500 9.8350 382.7500 10.1650 ;
        RECT 413.3500 9.8350 415.3500 10.1650 ;
        RECT 405.2000 9.8350 407.2000 10.1650 ;
        RECT 437.8000 9.8350 439.8000 10.1650 ;
        RECT 429.6500 9.8350 431.6500 10.1650 ;
        RECT 421.5000 9.8350 423.5000 10.1650 ;
        RECT 454.1000 9.8350 456.1000 10.1650 ;
        RECT 445.9500 9.8350 447.9500 10.1650 ;
        RECT 478.5500 9.8350 480.5500 10.1650 ;
        RECT 470.4000 9.8350 472.4000 10.1650 ;
        RECT 462.2500 9.8350 464.2500 10.1650 ;
        RECT 494.8500 9.8350 496.8500 10.1650 ;
        RECT 486.7000 9.8350 488.7000 10.1650 ;
        RECT 584.5000 9.8350 586.5000 10.1650 ;
        RECT 543.7500 9.8350 545.7500 10.1650 ;
        RECT 519.3000 9.8350 521.3000 10.1650 ;
        RECT 511.1500 9.8350 513.1500 10.1650 ;
        RECT 503.0000 9.8350 505.0000 10.1650 ;
        RECT 535.6000 9.8350 537.6000 10.1650 ;
        RECT 527.4500 9.8350 529.4500 10.1650 ;
        RECT 560.0500 9.8350 562.0500 10.1650 ;
        RECT 551.9000 9.8350 553.9000 10.1650 ;
        RECT 576.3500 9.8350 578.3500 10.1650 ;
        RECT 568.2000 9.8350 570.2000 10.1650 ;
        RECT 600.8000 9.8350 602.8000 10.1650 ;
        RECT 592.6500 9.8350 594.6500 10.1650 ;
        RECT 625.2500 9.8350 627.2500 10.1650 ;
        RECT 617.1000 9.8350 619.1000 10.1650 ;
        RECT 608.9500 9.8350 610.9500 10.1650 ;
        RECT 641.5500 9.8350 643.5500 10.1650 ;
        RECT 633.4000 9.8350 635.4000 10.1650 ;
        RECT 657.8500 9.8350 659.8500 10.1650 ;
        RECT 649.7000 9.8350 651.7000 10.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 670.0000 670.0000 ;
    LAYER M2 ;
      RECT 653.0500 669.3800 670.0000 670.0000 ;
      RECT 649.0500 669.3800 652.7500 670.0000 ;
      RECT 645.0500 669.3800 648.7500 670.0000 ;
      RECT 641.0500 669.3800 644.7500 670.0000 ;
      RECT 637.0500 669.3800 640.7500 670.0000 ;
      RECT 633.0500 669.3800 636.7500 670.0000 ;
      RECT 629.0500 669.3800 632.7500 670.0000 ;
      RECT 625.0500 669.3800 628.7500 670.0000 ;
      RECT 621.0500 669.3800 624.7500 670.0000 ;
      RECT 617.0500 669.3800 620.7500 670.0000 ;
      RECT 613.0500 669.3800 616.7500 670.0000 ;
      RECT 609.0500 669.3800 612.7500 670.0000 ;
      RECT 605.0500 669.3800 608.7500 670.0000 ;
      RECT 601.0500 669.3800 604.7500 670.0000 ;
      RECT 597.0500 669.3800 600.7500 670.0000 ;
      RECT 593.0500 669.3800 596.7500 670.0000 ;
      RECT 589.0500 669.3800 592.7500 670.0000 ;
      RECT 585.0500 669.3800 588.7500 670.0000 ;
      RECT 581.0500 669.3800 584.7500 670.0000 ;
      RECT 577.0500 669.3800 580.7500 670.0000 ;
      RECT 573.0500 669.3800 576.7500 670.0000 ;
      RECT 569.0500 669.3800 572.7500 670.0000 ;
      RECT 565.0500 669.3800 568.7500 670.0000 ;
      RECT 561.0500 669.3800 564.7500 670.0000 ;
      RECT 557.0500 669.3800 560.7500 670.0000 ;
      RECT 553.0500 669.3800 556.7500 670.0000 ;
      RECT 549.0500 669.3800 552.7500 670.0000 ;
      RECT 545.0500 669.3800 548.7500 670.0000 ;
      RECT 541.0500 669.3800 544.7500 670.0000 ;
      RECT 537.0500 669.3800 540.7500 670.0000 ;
      RECT 533.0500 669.3800 536.7500 670.0000 ;
      RECT 529.0500 669.3800 532.7500 670.0000 ;
      RECT 525.0500 669.3800 528.7500 670.0000 ;
      RECT 521.0500 669.3800 524.7500 670.0000 ;
      RECT 517.0500 669.3800 520.7500 670.0000 ;
      RECT 513.0500 669.3800 516.7500 670.0000 ;
      RECT 509.0500 669.3800 512.7500 670.0000 ;
      RECT 505.0500 669.3800 508.7500 670.0000 ;
      RECT 501.0500 669.3800 504.7500 670.0000 ;
      RECT 497.0500 669.3800 500.7500 670.0000 ;
      RECT 493.0500 669.3800 496.7500 670.0000 ;
      RECT 489.0500 669.3800 492.7500 670.0000 ;
      RECT 485.0500 669.3800 488.7500 670.0000 ;
      RECT 481.0500 669.3800 484.7500 670.0000 ;
      RECT 477.0500 669.3800 480.7500 670.0000 ;
      RECT 473.0500 669.3800 476.7500 670.0000 ;
      RECT 469.0500 669.3800 472.7500 670.0000 ;
      RECT 465.0500 669.3800 468.7500 670.0000 ;
      RECT 461.0500 669.3800 464.7500 670.0000 ;
      RECT 457.0500 669.3800 460.7500 670.0000 ;
      RECT 453.0500 669.3800 456.7500 670.0000 ;
      RECT 449.0500 669.3800 452.7500 670.0000 ;
      RECT 445.0500 669.3800 448.7500 670.0000 ;
      RECT 441.0500 669.3800 444.7500 670.0000 ;
      RECT 437.0500 669.3800 440.7500 670.0000 ;
      RECT 433.0500 669.3800 436.7500 670.0000 ;
      RECT 429.0500 669.3800 432.7500 670.0000 ;
      RECT 425.0500 669.3800 428.7500 670.0000 ;
      RECT 421.0500 669.3800 424.7500 670.0000 ;
      RECT 417.0500 669.3800 420.7500 670.0000 ;
      RECT 413.0500 669.3800 416.7500 670.0000 ;
      RECT 409.0500 669.3800 412.7500 670.0000 ;
      RECT 405.0500 669.3800 408.7500 670.0000 ;
      RECT 401.0500 669.3800 404.7500 670.0000 ;
      RECT 397.0500 669.3800 400.7500 670.0000 ;
      RECT 393.0500 669.3800 396.7500 670.0000 ;
      RECT 389.0500 669.3800 392.7500 670.0000 ;
      RECT 385.0500 669.3800 388.7500 670.0000 ;
      RECT 381.0500 669.3800 384.7500 670.0000 ;
      RECT 377.0500 669.3800 380.7500 670.0000 ;
      RECT 373.0500 669.3800 376.7500 670.0000 ;
      RECT 369.0500 669.3800 372.7500 670.0000 ;
      RECT 365.0500 669.3800 368.7500 670.0000 ;
      RECT 361.0500 669.3800 364.7500 670.0000 ;
      RECT 357.0500 669.3800 360.7500 670.0000 ;
      RECT 353.0500 669.3800 356.7500 670.0000 ;
      RECT 349.0500 669.3800 352.7500 670.0000 ;
      RECT 345.0500 669.3800 348.7500 670.0000 ;
      RECT 341.0500 669.3800 344.7500 670.0000 ;
      RECT 337.0500 669.3800 340.7500 670.0000 ;
      RECT 333.0500 669.3800 336.7500 670.0000 ;
      RECT 329.0500 669.3800 332.7500 670.0000 ;
      RECT 325.0500 669.3800 328.7500 670.0000 ;
      RECT 321.0500 669.3800 324.7500 670.0000 ;
      RECT 317.0500 669.3800 320.7500 670.0000 ;
      RECT 313.0500 669.3800 316.7500 670.0000 ;
      RECT 309.0500 669.3800 312.7500 670.0000 ;
      RECT 305.0500 669.3800 308.7500 670.0000 ;
      RECT 301.0500 669.3800 304.7500 670.0000 ;
      RECT 297.0500 669.3800 300.7500 670.0000 ;
      RECT 293.0500 669.3800 296.7500 670.0000 ;
      RECT 289.0500 669.3800 292.7500 670.0000 ;
      RECT 285.0500 669.3800 288.7500 670.0000 ;
      RECT 281.0500 669.3800 284.7500 670.0000 ;
      RECT 277.0500 669.3800 280.7500 670.0000 ;
      RECT 273.0500 669.3800 276.7500 670.0000 ;
      RECT 269.0500 669.3800 272.7500 670.0000 ;
      RECT 265.0500 669.3800 268.7500 670.0000 ;
      RECT 261.0500 669.3800 264.7500 670.0000 ;
      RECT 257.0500 669.3800 260.7500 670.0000 ;
      RECT 253.0500 669.3800 256.7500 670.0000 ;
      RECT 249.0500 669.3800 252.7500 670.0000 ;
      RECT 245.0500 669.3800 248.7500 670.0000 ;
      RECT 241.0500 669.3800 244.7500 670.0000 ;
      RECT 237.0500 669.3800 240.7500 670.0000 ;
      RECT 233.0500 669.3800 236.7500 670.0000 ;
      RECT 229.0500 669.3800 232.7500 670.0000 ;
      RECT 225.0500 669.3800 228.7500 670.0000 ;
      RECT 221.0500 669.3800 224.7500 670.0000 ;
      RECT 217.0500 669.3800 220.7500 670.0000 ;
      RECT 213.0500 669.3800 216.7500 670.0000 ;
      RECT 209.0500 669.3800 212.7500 670.0000 ;
      RECT 205.0500 669.3800 208.7500 670.0000 ;
      RECT 201.0500 669.3800 204.7500 670.0000 ;
      RECT 197.0500 669.3800 200.7500 670.0000 ;
      RECT 193.0500 669.3800 196.7500 670.0000 ;
      RECT 189.0500 669.3800 192.7500 670.0000 ;
      RECT 185.0500 669.3800 188.7500 670.0000 ;
      RECT 181.0500 669.3800 184.7500 670.0000 ;
      RECT 177.0500 669.3800 180.7500 670.0000 ;
      RECT 173.0500 669.3800 176.7500 670.0000 ;
      RECT 169.0500 669.3800 172.7500 670.0000 ;
      RECT 165.0500 669.3800 168.7500 670.0000 ;
      RECT 161.0500 669.3800 164.7500 670.0000 ;
      RECT 157.0500 669.3800 160.7500 670.0000 ;
      RECT 153.0500 669.3800 156.7500 670.0000 ;
      RECT 149.0500 669.3800 152.7500 670.0000 ;
      RECT 145.0500 669.3800 148.7500 670.0000 ;
      RECT 141.0500 669.3800 144.7500 670.0000 ;
      RECT 137.0500 669.3800 140.7500 670.0000 ;
      RECT 133.0500 669.3800 136.7500 670.0000 ;
      RECT 129.0500 669.3800 132.7500 670.0000 ;
      RECT 125.0500 669.3800 128.7500 670.0000 ;
      RECT 121.0500 669.3800 124.7500 670.0000 ;
      RECT 117.0500 669.3800 120.7500 670.0000 ;
      RECT 113.0500 669.3800 116.7500 670.0000 ;
      RECT 109.0500 669.3800 112.7500 670.0000 ;
      RECT 105.0500 669.3800 108.7500 670.0000 ;
      RECT 101.0500 669.3800 104.7500 670.0000 ;
      RECT 97.0500 669.3800 100.7500 670.0000 ;
      RECT 93.0500 669.3800 96.7500 670.0000 ;
      RECT 89.0500 669.3800 92.7500 670.0000 ;
      RECT 85.0500 669.3800 88.7500 670.0000 ;
      RECT 81.0500 669.3800 84.7500 670.0000 ;
      RECT 77.0500 669.3800 80.7500 670.0000 ;
      RECT 73.0500 669.3800 76.7500 670.0000 ;
      RECT 69.0500 669.3800 72.7500 670.0000 ;
      RECT 65.0500 669.3800 68.7500 670.0000 ;
      RECT 61.0500 669.3800 64.7500 670.0000 ;
      RECT 57.0500 669.3800 60.7500 670.0000 ;
      RECT 53.0500 669.3800 56.7500 670.0000 ;
      RECT 49.0500 669.3800 52.7500 670.0000 ;
      RECT 45.0500 669.3800 48.7500 670.0000 ;
      RECT 41.0500 669.3800 44.7500 670.0000 ;
      RECT 37.0500 669.3800 40.7500 670.0000 ;
      RECT 33.0500 669.3800 36.7500 670.0000 ;
      RECT 29.0500 669.3800 32.7500 670.0000 ;
      RECT 25.0500 669.3800 28.7500 670.0000 ;
      RECT 21.0500 669.3800 24.7500 670.0000 ;
      RECT 17.0500 669.3800 20.7500 670.0000 ;
      RECT 0.0000 669.3800 16.7500 670.0000 ;
      RECT 0.0000 0.6200 670.0000 669.3800 ;
      RECT 653.0500 0.0000 670.0000 0.6200 ;
      RECT 649.0500 0.0000 652.7500 0.6200 ;
      RECT 645.0500 0.0000 648.7500 0.6200 ;
      RECT 641.0500 0.0000 644.7500 0.6200 ;
      RECT 637.0500 0.0000 640.7500 0.6200 ;
      RECT 633.0500 0.0000 636.7500 0.6200 ;
      RECT 629.0500 0.0000 632.7500 0.6200 ;
      RECT 625.0500 0.0000 628.7500 0.6200 ;
      RECT 621.0500 0.0000 624.7500 0.6200 ;
      RECT 617.0500 0.0000 620.7500 0.6200 ;
      RECT 613.0500 0.0000 616.7500 0.6200 ;
      RECT 609.0500 0.0000 612.7500 0.6200 ;
      RECT 605.0500 0.0000 608.7500 0.6200 ;
      RECT 601.0500 0.0000 604.7500 0.6200 ;
      RECT 597.0500 0.0000 600.7500 0.6200 ;
      RECT 593.0500 0.0000 596.7500 0.6200 ;
      RECT 589.0500 0.0000 592.7500 0.6200 ;
      RECT 585.0500 0.0000 588.7500 0.6200 ;
      RECT 581.0500 0.0000 584.7500 0.6200 ;
      RECT 577.0500 0.0000 580.7500 0.6200 ;
      RECT 573.0500 0.0000 576.7500 0.6200 ;
      RECT 569.0500 0.0000 572.7500 0.6200 ;
      RECT 565.0500 0.0000 568.7500 0.6200 ;
      RECT 561.0500 0.0000 564.7500 0.6200 ;
      RECT 557.0500 0.0000 560.7500 0.6200 ;
      RECT 553.0500 0.0000 556.7500 0.6200 ;
      RECT 549.0500 0.0000 552.7500 0.6200 ;
      RECT 545.0500 0.0000 548.7500 0.6200 ;
      RECT 541.0500 0.0000 544.7500 0.6200 ;
      RECT 537.0500 0.0000 540.7500 0.6200 ;
      RECT 533.0500 0.0000 536.7500 0.6200 ;
      RECT 529.0500 0.0000 532.7500 0.6200 ;
      RECT 525.0500 0.0000 528.7500 0.6200 ;
      RECT 521.0500 0.0000 524.7500 0.6200 ;
      RECT 517.0500 0.0000 520.7500 0.6200 ;
      RECT 513.0500 0.0000 516.7500 0.6200 ;
      RECT 509.0500 0.0000 512.7500 0.6200 ;
      RECT 505.0500 0.0000 508.7500 0.6200 ;
      RECT 501.0500 0.0000 504.7500 0.6200 ;
      RECT 497.0500 0.0000 500.7500 0.6200 ;
      RECT 493.0500 0.0000 496.7500 0.6200 ;
      RECT 489.0500 0.0000 492.7500 0.6200 ;
      RECT 485.0500 0.0000 488.7500 0.6200 ;
      RECT 481.0500 0.0000 484.7500 0.6200 ;
      RECT 477.0500 0.0000 480.7500 0.6200 ;
      RECT 473.0500 0.0000 476.7500 0.6200 ;
      RECT 469.0500 0.0000 472.7500 0.6200 ;
      RECT 465.0500 0.0000 468.7500 0.6200 ;
      RECT 461.0500 0.0000 464.7500 0.6200 ;
      RECT 457.0500 0.0000 460.7500 0.6200 ;
      RECT 453.0500 0.0000 456.7500 0.6200 ;
      RECT 449.0500 0.0000 452.7500 0.6200 ;
      RECT 445.0500 0.0000 448.7500 0.6200 ;
      RECT 441.0500 0.0000 444.7500 0.6200 ;
      RECT 437.0500 0.0000 440.7500 0.6200 ;
      RECT 433.0500 0.0000 436.7500 0.6200 ;
      RECT 429.0500 0.0000 432.7500 0.6200 ;
      RECT 425.0500 0.0000 428.7500 0.6200 ;
      RECT 421.0500 0.0000 424.7500 0.6200 ;
      RECT 417.0500 0.0000 420.7500 0.6200 ;
      RECT 413.0500 0.0000 416.7500 0.6200 ;
      RECT 409.0500 0.0000 412.7500 0.6200 ;
      RECT 405.0500 0.0000 408.7500 0.6200 ;
      RECT 401.0500 0.0000 404.7500 0.6200 ;
      RECT 397.0500 0.0000 400.7500 0.6200 ;
      RECT 393.0500 0.0000 396.7500 0.6200 ;
      RECT 389.0500 0.0000 392.7500 0.6200 ;
      RECT 385.0500 0.0000 388.7500 0.6200 ;
      RECT 381.0500 0.0000 384.7500 0.6200 ;
      RECT 377.0500 0.0000 380.7500 0.6200 ;
      RECT 373.0500 0.0000 376.7500 0.6200 ;
      RECT 369.0500 0.0000 372.7500 0.6200 ;
      RECT 365.0500 0.0000 368.7500 0.6200 ;
      RECT 361.0500 0.0000 364.7500 0.6200 ;
      RECT 357.0500 0.0000 360.7500 0.6200 ;
      RECT 353.0500 0.0000 356.7500 0.6200 ;
      RECT 349.0500 0.0000 352.7500 0.6200 ;
      RECT 345.0500 0.0000 348.7500 0.6200 ;
      RECT 341.0500 0.0000 344.7500 0.6200 ;
      RECT 337.0500 0.0000 340.7500 0.6200 ;
      RECT 333.0500 0.0000 336.7500 0.6200 ;
      RECT 329.0500 0.0000 332.7500 0.6200 ;
      RECT 325.0500 0.0000 328.7500 0.6200 ;
      RECT 321.0500 0.0000 324.7500 0.6200 ;
      RECT 317.0500 0.0000 320.7500 0.6200 ;
      RECT 313.0500 0.0000 316.7500 0.6200 ;
      RECT 309.0500 0.0000 312.7500 0.6200 ;
      RECT 305.0500 0.0000 308.7500 0.6200 ;
      RECT 301.0500 0.0000 304.7500 0.6200 ;
      RECT 297.0500 0.0000 300.7500 0.6200 ;
      RECT 293.0500 0.0000 296.7500 0.6200 ;
      RECT 289.0500 0.0000 292.7500 0.6200 ;
      RECT 285.0500 0.0000 288.7500 0.6200 ;
      RECT 281.0500 0.0000 284.7500 0.6200 ;
      RECT 277.0500 0.0000 280.7500 0.6200 ;
      RECT 273.0500 0.0000 276.7500 0.6200 ;
      RECT 269.0500 0.0000 272.7500 0.6200 ;
      RECT 265.0500 0.0000 268.7500 0.6200 ;
      RECT 261.0500 0.0000 264.7500 0.6200 ;
      RECT 257.0500 0.0000 260.7500 0.6200 ;
      RECT 253.0500 0.0000 256.7500 0.6200 ;
      RECT 249.0500 0.0000 252.7500 0.6200 ;
      RECT 245.0500 0.0000 248.7500 0.6200 ;
      RECT 241.0500 0.0000 244.7500 0.6200 ;
      RECT 237.0500 0.0000 240.7500 0.6200 ;
      RECT 233.0500 0.0000 236.7500 0.6200 ;
      RECT 229.0500 0.0000 232.7500 0.6200 ;
      RECT 225.0500 0.0000 228.7500 0.6200 ;
      RECT 221.0500 0.0000 224.7500 0.6200 ;
      RECT 217.0500 0.0000 220.7500 0.6200 ;
      RECT 213.0500 0.0000 216.7500 0.6200 ;
      RECT 209.0500 0.0000 212.7500 0.6200 ;
      RECT 205.0500 0.0000 208.7500 0.6200 ;
      RECT 201.0500 0.0000 204.7500 0.6200 ;
      RECT 197.0500 0.0000 200.7500 0.6200 ;
      RECT 193.0500 0.0000 196.7500 0.6200 ;
      RECT 189.0500 0.0000 192.7500 0.6200 ;
      RECT 185.0500 0.0000 188.7500 0.6200 ;
      RECT 181.0500 0.0000 184.7500 0.6200 ;
      RECT 177.0500 0.0000 180.7500 0.6200 ;
      RECT 173.0500 0.0000 176.7500 0.6200 ;
      RECT 169.0500 0.0000 172.7500 0.6200 ;
      RECT 165.0500 0.0000 168.7500 0.6200 ;
      RECT 161.0500 0.0000 164.7500 0.6200 ;
      RECT 157.0500 0.0000 160.7500 0.6200 ;
      RECT 153.0500 0.0000 156.7500 0.6200 ;
      RECT 149.0500 0.0000 152.7500 0.6200 ;
      RECT 145.0500 0.0000 148.7500 0.6200 ;
      RECT 141.0500 0.0000 144.7500 0.6200 ;
      RECT 137.0500 0.0000 140.7500 0.6200 ;
      RECT 133.0500 0.0000 136.7500 0.6200 ;
      RECT 129.0500 0.0000 132.7500 0.6200 ;
      RECT 125.0500 0.0000 128.7500 0.6200 ;
      RECT 121.0500 0.0000 124.7500 0.6200 ;
      RECT 117.0500 0.0000 120.7500 0.6200 ;
      RECT 113.0500 0.0000 116.7500 0.6200 ;
      RECT 109.0500 0.0000 112.7500 0.6200 ;
      RECT 105.0500 0.0000 108.7500 0.6200 ;
      RECT 101.0500 0.0000 104.7500 0.6200 ;
      RECT 97.0500 0.0000 100.7500 0.6200 ;
      RECT 93.0500 0.0000 96.7500 0.6200 ;
      RECT 89.0500 0.0000 92.7500 0.6200 ;
      RECT 85.0500 0.0000 88.7500 0.6200 ;
      RECT 81.0500 0.0000 84.7500 0.6200 ;
      RECT 77.0500 0.0000 80.7500 0.6200 ;
      RECT 73.0500 0.0000 76.7500 0.6200 ;
      RECT 69.0500 0.0000 72.7500 0.6200 ;
      RECT 65.0500 0.0000 68.7500 0.6200 ;
      RECT 61.0500 0.0000 64.7500 0.6200 ;
      RECT 57.0500 0.0000 60.7500 0.6200 ;
      RECT 53.0500 0.0000 56.7500 0.6200 ;
      RECT 49.0500 0.0000 52.7500 0.6200 ;
      RECT 45.0500 0.0000 48.7500 0.6200 ;
      RECT 41.0500 0.0000 44.7500 0.6200 ;
      RECT 37.0500 0.0000 40.7500 0.6200 ;
      RECT 33.0500 0.0000 36.7500 0.6200 ;
      RECT 29.0500 0.0000 32.7500 0.6200 ;
      RECT 25.0500 0.0000 28.7500 0.6200 ;
      RECT 21.0500 0.0000 24.7500 0.6200 ;
      RECT 17.0500 0.0000 20.7500 0.6200 ;
      RECT 0.0000 0.0000 16.7500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 346.9500 670.0000 670.0000 ;
      RECT 0.6200 346.6500 670.0000 346.9500 ;
      RECT 0.0000 342.9500 670.0000 346.6500 ;
      RECT 0.6200 342.6500 670.0000 342.9500 ;
      RECT 0.0000 338.9500 670.0000 342.6500 ;
      RECT 0.6200 338.6500 670.0000 338.9500 ;
      RECT 0.0000 334.9500 670.0000 338.6500 ;
      RECT 0.6200 334.6500 670.0000 334.9500 ;
      RECT 0.0000 330.9500 670.0000 334.6500 ;
      RECT 0.6200 330.6500 670.0000 330.9500 ;
      RECT 0.0000 326.9500 670.0000 330.6500 ;
      RECT 0.6200 326.6500 670.0000 326.9500 ;
      RECT 0.0000 322.9500 670.0000 326.6500 ;
      RECT 0.6200 322.6500 670.0000 322.9500 ;
      RECT 0.0000 0.0000 670.0000 322.6500 ;
    LAYER M4 ;
      RECT 0.0000 660.5000 670.0000 670.0000 ;
      RECT 656.3500 9.5000 657.3500 660.5000 ;
      RECT 652.2000 9.5000 653.3500 660.5000 ;
      RECT 648.2000 9.5000 649.2000 660.5000 ;
      RECT 644.0500 9.5000 645.2000 660.5000 ;
      RECT 640.0500 9.5000 641.0500 660.5000 ;
      RECT 635.9000 9.5000 637.0500 660.5000 ;
      RECT 631.9000 9.5000 632.9000 660.5000 ;
      RECT 627.7500 9.5000 628.9000 660.5000 ;
      RECT 623.7500 9.5000 624.7500 660.5000 ;
      RECT 619.6000 9.5000 620.7500 660.5000 ;
      RECT 615.6000 9.5000 616.6000 660.5000 ;
      RECT 611.4500 9.5000 612.6000 660.5000 ;
      RECT 607.4500 9.5000 608.4500 660.5000 ;
      RECT 603.3000 9.5000 604.4500 660.5000 ;
      RECT 599.3000 9.5000 600.3000 660.5000 ;
      RECT 595.1500 9.5000 596.3000 660.5000 ;
      RECT 591.1500 9.5000 592.1500 660.5000 ;
      RECT 587.0000 9.5000 588.1500 660.5000 ;
      RECT 583.0000 9.5000 584.0000 660.5000 ;
      RECT 578.8500 9.5000 580.0000 660.5000 ;
      RECT 574.8500 9.5000 575.8500 660.5000 ;
      RECT 570.7000 9.5000 571.8500 660.5000 ;
      RECT 566.7000 9.5000 567.7000 660.5000 ;
      RECT 562.5500 9.5000 563.7000 660.5000 ;
      RECT 558.5500 9.5000 559.5500 660.5000 ;
      RECT 554.4000 9.5000 555.5500 660.5000 ;
      RECT 550.4000 9.5000 551.4000 660.5000 ;
      RECT 546.2500 9.5000 547.4000 660.5000 ;
      RECT 542.2500 9.5000 543.2500 660.5000 ;
      RECT 538.1000 9.5000 539.2500 660.5000 ;
      RECT 534.1000 9.5000 535.1000 660.5000 ;
      RECT 529.9500 9.5000 531.1000 660.5000 ;
      RECT 525.9500 9.5000 526.9500 660.5000 ;
      RECT 521.8000 9.5000 522.9500 660.5000 ;
      RECT 517.8000 9.5000 518.8000 660.5000 ;
      RECT 513.6500 9.5000 514.8000 660.5000 ;
      RECT 509.6500 9.5000 510.6500 660.5000 ;
      RECT 505.5000 9.5000 506.6500 660.5000 ;
      RECT 501.5000 9.5000 502.5000 660.5000 ;
      RECT 497.3500 9.5000 498.5000 660.5000 ;
      RECT 493.3500 9.5000 494.3500 660.5000 ;
      RECT 489.2000 9.5000 490.3500 660.5000 ;
      RECT 485.2000 9.5000 486.2000 660.5000 ;
      RECT 481.0500 9.5000 482.2000 660.5000 ;
      RECT 477.0500 9.5000 478.0500 660.5000 ;
      RECT 472.9000 9.5000 474.0500 660.5000 ;
      RECT 468.9000 9.5000 469.9000 660.5000 ;
      RECT 464.7500 9.5000 465.9000 660.5000 ;
      RECT 460.7500 9.5000 461.7500 660.5000 ;
      RECT 456.6000 9.5000 457.7500 660.5000 ;
      RECT 452.6000 9.5000 453.6000 660.5000 ;
      RECT 448.4500 9.5000 449.6000 660.5000 ;
      RECT 444.4500 9.5000 445.4500 660.5000 ;
      RECT 440.3000 9.5000 441.4500 660.5000 ;
      RECT 436.3000 9.5000 437.3000 660.5000 ;
      RECT 432.1500 9.5000 433.3000 660.5000 ;
      RECT 428.1500 9.5000 429.1500 660.5000 ;
      RECT 424.0000 9.5000 425.1500 660.5000 ;
      RECT 420.0000 9.5000 421.0000 660.5000 ;
      RECT 415.8500 9.5000 417.0000 660.5000 ;
      RECT 411.8500 9.5000 412.8500 660.5000 ;
      RECT 407.7000 9.5000 408.8500 660.5000 ;
      RECT 403.7000 9.5000 404.7000 660.5000 ;
      RECT 399.5500 9.5000 400.7000 660.5000 ;
      RECT 395.5500 9.5000 396.5500 660.5000 ;
      RECT 391.4000 9.5000 392.5500 660.5000 ;
      RECT 387.4000 9.5000 388.4000 660.5000 ;
      RECT 383.2500 9.5000 384.4000 660.5000 ;
      RECT 379.2500 9.5000 380.2500 660.5000 ;
      RECT 375.1000 9.5000 376.2500 660.5000 ;
      RECT 371.1000 9.5000 372.1000 660.5000 ;
      RECT 366.9500 9.5000 368.1000 660.5000 ;
      RECT 362.9500 9.5000 363.9500 660.5000 ;
      RECT 358.8000 9.5000 359.9500 660.5000 ;
      RECT 354.8000 9.5000 355.8000 660.5000 ;
      RECT 350.6500 9.5000 351.8000 660.5000 ;
      RECT 346.6500 9.5000 347.6500 660.5000 ;
      RECT 342.5000 9.5000 343.6500 660.5000 ;
      RECT 338.5000 9.5000 339.5000 660.5000 ;
      RECT 334.3500 9.5000 335.5000 660.5000 ;
      RECT 330.3500 9.5000 331.3500 660.5000 ;
      RECT 326.2000 9.5000 327.3500 660.5000 ;
      RECT 322.2000 9.5000 323.2000 660.5000 ;
      RECT 318.0500 9.5000 319.2000 660.5000 ;
      RECT 314.0500 9.5000 315.0500 660.5000 ;
      RECT 309.9000 9.5000 311.0500 660.5000 ;
      RECT 305.9000 9.5000 306.9000 660.5000 ;
      RECT 301.7500 9.5000 302.9000 660.5000 ;
      RECT 297.7500 9.5000 298.7500 660.5000 ;
      RECT 293.6000 9.5000 294.7500 660.5000 ;
      RECT 289.6000 9.5000 290.6000 660.5000 ;
      RECT 285.4500 9.5000 286.6000 660.5000 ;
      RECT 281.4500 9.5000 282.4500 660.5000 ;
      RECT 277.3000 9.5000 278.4500 660.5000 ;
      RECT 273.3000 9.5000 274.3000 660.5000 ;
      RECT 269.1500 9.5000 270.3000 660.5000 ;
      RECT 265.1500 9.5000 266.1500 660.5000 ;
      RECT 261.0000 9.5000 262.1500 660.5000 ;
      RECT 257.0000 9.5000 258.0000 660.5000 ;
      RECT 252.8500 9.5000 254.0000 660.5000 ;
      RECT 248.8500 9.5000 249.8500 660.5000 ;
      RECT 244.7000 9.5000 245.8500 660.5000 ;
      RECT 240.7000 9.5000 241.7000 660.5000 ;
      RECT 236.5500 9.5000 237.7000 660.5000 ;
      RECT 232.5500 9.5000 233.5500 660.5000 ;
      RECT 228.4000 9.5000 229.5500 660.5000 ;
      RECT 224.4000 9.5000 225.4000 660.5000 ;
      RECT 220.2500 9.5000 221.4000 660.5000 ;
      RECT 216.2500 9.5000 217.2500 660.5000 ;
      RECT 212.1000 9.5000 213.2500 660.5000 ;
      RECT 208.1000 9.5000 209.1000 660.5000 ;
      RECT 203.9500 9.5000 205.1000 660.5000 ;
      RECT 199.9500 9.5000 200.9500 660.5000 ;
      RECT 195.8000 9.5000 196.9500 660.5000 ;
      RECT 191.8000 9.5000 192.8000 660.5000 ;
      RECT 187.6500 9.5000 188.8000 660.5000 ;
      RECT 183.6500 9.5000 184.6500 660.5000 ;
      RECT 179.5000 9.5000 180.6500 660.5000 ;
      RECT 175.5000 9.5000 176.5000 660.5000 ;
      RECT 171.3500 9.5000 172.5000 660.5000 ;
      RECT 167.3500 9.5000 168.3500 660.5000 ;
      RECT 163.2000 9.5000 164.3500 660.5000 ;
      RECT 159.2000 9.5000 160.2000 660.5000 ;
      RECT 155.0500 9.5000 156.2000 660.5000 ;
      RECT 151.0500 9.5000 152.0500 660.5000 ;
      RECT 146.9000 9.5000 148.0500 660.5000 ;
      RECT 142.9000 9.5000 143.9000 660.5000 ;
      RECT 138.7500 9.5000 139.9000 660.5000 ;
      RECT 134.7500 9.5000 135.7500 660.5000 ;
      RECT 130.6000 9.5000 131.7500 660.5000 ;
      RECT 126.6000 9.5000 127.6000 660.5000 ;
      RECT 122.4500 9.5000 123.6000 660.5000 ;
      RECT 118.4500 9.5000 119.4500 660.5000 ;
      RECT 114.3000 9.5000 115.4500 660.5000 ;
      RECT 110.3000 9.5000 111.3000 660.5000 ;
      RECT 106.1500 9.5000 107.3000 660.5000 ;
      RECT 102.1500 9.5000 103.1500 660.5000 ;
      RECT 98.0000 9.5000 99.1500 660.5000 ;
      RECT 94.0000 9.5000 95.0000 660.5000 ;
      RECT 89.8500 9.5000 91.0000 660.5000 ;
      RECT 85.8500 9.5000 86.8500 660.5000 ;
      RECT 81.7000 9.5000 82.8500 660.5000 ;
      RECT 77.7000 9.5000 78.7000 660.5000 ;
      RECT 73.5500 9.5000 74.7000 660.5000 ;
      RECT 69.5500 9.5000 70.5500 660.5000 ;
      RECT 65.4000 9.5000 66.5500 660.5000 ;
      RECT 61.4000 9.5000 62.4000 660.5000 ;
      RECT 57.2500 9.5000 58.4000 660.5000 ;
      RECT 53.2500 9.5000 54.2500 660.5000 ;
      RECT 49.1000 9.5000 50.2500 660.5000 ;
      RECT 45.1000 9.5000 46.1000 660.5000 ;
      RECT 40.9500 9.5000 42.1000 660.5000 ;
      RECT 36.9500 9.5000 37.9500 660.5000 ;
      RECT 32.8000 9.5000 33.9500 660.5000 ;
      RECT 28.8000 9.5000 29.8000 660.5000 ;
      RECT 24.6500 9.5000 25.8000 660.5000 ;
      RECT 20.6500 9.5000 21.6500 660.5000 ;
      RECT 16.5000 9.5000 17.6500 660.5000 ;
      RECT 12.5000 9.5000 13.5000 660.5000 ;
      RECT 0.0000 9.5000 9.5000 660.5000 ;
      RECT 660.3500 9.3350 670.0000 660.5000 ;
      RECT 652.2000 9.3350 657.3500 9.5000 ;
      RECT 644.0500 9.3350 649.2000 9.5000 ;
      RECT 635.9000 9.3350 641.0500 9.5000 ;
      RECT 627.7500 9.3350 632.9000 9.5000 ;
      RECT 619.6000 9.3350 624.7500 9.5000 ;
      RECT 611.4500 9.3350 616.6000 9.5000 ;
      RECT 603.3000 9.3350 608.4500 9.5000 ;
      RECT 595.1500 9.3350 600.3000 9.5000 ;
      RECT 587.0000 9.3350 592.1500 9.5000 ;
      RECT 578.8500 9.3350 584.0000 9.5000 ;
      RECT 570.7000 9.3350 575.8500 9.5000 ;
      RECT 562.5500 9.3350 567.7000 9.5000 ;
      RECT 554.4000 9.3350 559.5500 9.5000 ;
      RECT 546.2500 9.3350 551.4000 9.5000 ;
      RECT 538.1000 9.3350 543.2500 9.5000 ;
      RECT 529.9500 9.3350 535.1000 9.5000 ;
      RECT 521.8000 9.3350 526.9500 9.5000 ;
      RECT 513.6500 9.3350 518.8000 9.5000 ;
      RECT 505.5000 9.3350 510.6500 9.5000 ;
      RECT 497.3500 9.3350 502.5000 9.5000 ;
      RECT 489.2000 9.3350 494.3500 9.5000 ;
      RECT 481.0500 9.3350 486.2000 9.5000 ;
      RECT 472.9000 9.3350 478.0500 9.5000 ;
      RECT 464.7500 9.3350 469.9000 9.5000 ;
      RECT 456.6000 9.3350 461.7500 9.5000 ;
      RECT 448.4500 9.3350 453.6000 9.5000 ;
      RECT 440.3000 9.3350 445.4500 9.5000 ;
      RECT 432.1500 9.3350 437.3000 9.5000 ;
      RECT 424.0000 9.3350 429.1500 9.5000 ;
      RECT 415.8500 9.3350 421.0000 9.5000 ;
      RECT 407.7000 9.3350 412.8500 9.5000 ;
      RECT 399.5500 9.3350 404.7000 9.5000 ;
      RECT 391.4000 9.3350 396.5500 9.5000 ;
      RECT 383.2500 9.3350 388.4000 9.5000 ;
      RECT 375.1000 9.3350 380.2500 9.5000 ;
      RECT 366.9500 9.3350 372.1000 9.5000 ;
      RECT 358.8000 9.3350 363.9500 9.5000 ;
      RECT 350.6500 9.3350 355.8000 9.5000 ;
      RECT 342.5000 9.3350 347.6500 9.5000 ;
      RECT 334.3500 9.3350 339.5000 9.5000 ;
      RECT 326.2000 9.3350 331.3500 9.5000 ;
      RECT 318.0500 9.3350 323.2000 9.5000 ;
      RECT 309.9000 9.3350 315.0500 9.5000 ;
      RECT 301.7500 9.3350 306.9000 9.5000 ;
      RECT 293.6000 9.3350 298.7500 9.5000 ;
      RECT 285.4500 9.3350 290.6000 9.5000 ;
      RECT 277.3000 9.3350 282.4500 9.5000 ;
      RECT 269.1500 9.3350 274.3000 9.5000 ;
      RECT 261.0000 9.3350 266.1500 9.5000 ;
      RECT 252.8500 9.3350 258.0000 9.5000 ;
      RECT 244.7000 9.3350 249.8500 9.5000 ;
      RECT 236.5500 9.3350 241.7000 9.5000 ;
      RECT 228.4000 9.3350 233.5500 9.5000 ;
      RECT 220.2500 9.3350 225.4000 9.5000 ;
      RECT 212.1000 9.3350 217.2500 9.5000 ;
      RECT 203.9500 9.3350 209.1000 9.5000 ;
      RECT 195.8000 9.3350 200.9500 9.5000 ;
      RECT 187.6500 9.3350 192.8000 9.5000 ;
      RECT 179.5000 9.3350 184.6500 9.5000 ;
      RECT 171.3500 9.3350 176.5000 9.5000 ;
      RECT 163.2000 9.3350 168.3500 9.5000 ;
      RECT 155.0500 9.3350 160.2000 9.5000 ;
      RECT 146.9000 9.3350 152.0500 9.5000 ;
      RECT 138.7500 9.3350 143.9000 9.5000 ;
      RECT 130.6000 9.3350 135.7500 9.5000 ;
      RECT 122.4500 9.3350 127.6000 9.5000 ;
      RECT 114.3000 9.3350 119.4500 9.5000 ;
      RECT 106.1500 9.3350 111.3000 9.5000 ;
      RECT 98.0000 9.3350 103.1500 9.5000 ;
      RECT 89.8500 9.3350 95.0000 9.5000 ;
      RECT 81.7000 9.3350 86.8500 9.5000 ;
      RECT 73.5500 9.3350 78.7000 9.5000 ;
      RECT 65.4000 9.3350 70.5500 9.5000 ;
      RECT 57.2500 9.3350 62.4000 9.5000 ;
      RECT 49.1000 9.3350 54.2500 9.5000 ;
      RECT 40.9500 9.3350 46.1000 9.5000 ;
      RECT 32.8000 9.3350 37.9500 9.5000 ;
      RECT 24.6500 9.3350 29.8000 9.5000 ;
      RECT 16.5000 9.3350 21.6500 9.5000 ;
      RECT 0.0000 9.3350 13.5000 9.5000 ;
      RECT 0.0000 0.0000 670.0000 9.3350 ;
  END
END sram_w16_160b

END LIBRARY
