##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 10:54:32 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 1420.0000 BY 2820.0000 ;
  FOREIGN fullchip 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 418.0500 0.0000 418.1500 0.5200 ;
    END
  END clk
  PIN mem_in_core0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 498.0500 0.0000 498.1500 0.5200 ;
    END
  END mem_in_core0[63]
  PIN mem_in_core0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 502.0500 0.0000 502.1500 0.5200 ;
    END
  END mem_in_core0[62]
  PIN mem_in_core0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 506.0500 0.0000 506.1500 0.5200 ;
    END
  END mem_in_core0[61]
  PIN mem_in_core0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 510.0500 0.0000 510.1500 0.5200 ;
    END
  END mem_in_core0[60]
  PIN mem_in_core0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 514.0500 0.0000 514.1500 0.5200 ;
    END
  END mem_in_core0[59]
  PIN mem_in_core0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 518.0500 0.0000 518.1500 0.5200 ;
    END
  END mem_in_core0[58]
  PIN mem_in_core0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 522.0500 0.0000 522.1500 0.5200 ;
    END
  END mem_in_core0[57]
  PIN mem_in_core0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 526.0500 0.0000 526.1500 0.5200 ;
    END
  END mem_in_core0[56]
  PIN mem_in_core0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 530.0500 0.0000 530.1500 0.5200 ;
    END
  END mem_in_core0[55]
  PIN mem_in_core0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 534.0500 0.0000 534.1500 0.5200 ;
    END
  END mem_in_core0[54]
  PIN mem_in_core0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 538.0500 0.0000 538.1500 0.5200 ;
    END
  END mem_in_core0[53]
  PIN mem_in_core0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 542.0500 0.0000 542.1500 0.5200 ;
    END
  END mem_in_core0[52]
  PIN mem_in_core0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 546.0500 0.0000 546.1500 0.5200 ;
    END
  END mem_in_core0[51]
  PIN mem_in_core0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 550.0500 0.0000 550.1500 0.5200 ;
    END
  END mem_in_core0[50]
  PIN mem_in_core0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 554.0500 0.0000 554.1500 0.5200 ;
    END
  END mem_in_core0[49]
  PIN mem_in_core0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 558.0500 0.0000 558.1500 0.5200 ;
    END
  END mem_in_core0[48]
  PIN mem_in_core0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 562.0500 0.0000 562.1500 0.5200 ;
    END
  END mem_in_core0[47]
  PIN mem_in_core0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 566.0500 0.0000 566.1500 0.5200 ;
    END
  END mem_in_core0[46]
  PIN mem_in_core0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 570.0500 0.0000 570.1500 0.5200 ;
    END
  END mem_in_core0[45]
  PIN mem_in_core0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 574.0500 0.0000 574.1500 0.5200 ;
    END
  END mem_in_core0[44]
  PIN mem_in_core0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 578.0500 0.0000 578.1500 0.5200 ;
    END
  END mem_in_core0[43]
  PIN mem_in_core0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 582.0500 0.0000 582.1500 0.5200 ;
    END
  END mem_in_core0[42]
  PIN mem_in_core0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 586.0500 0.0000 586.1500 0.5200 ;
    END
  END mem_in_core0[41]
  PIN mem_in_core0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 590.0500 0.0000 590.1500 0.5200 ;
    END
  END mem_in_core0[40]
  PIN mem_in_core0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 594.0500 0.0000 594.1500 0.5200 ;
    END
  END mem_in_core0[39]
  PIN mem_in_core0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 598.0500 0.0000 598.1500 0.5200 ;
    END
  END mem_in_core0[38]
  PIN mem_in_core0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 602.0500 0.0000 602.1500 0.5200 ;
    END
  END mem_in_core0[37]
  PIN mem_in_core0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 606.0500 0.0000 606.1500 0.5200 ;
    END
  END mem_in_core0[36]
  PIN mem_in_core0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 610.0500 0.0000 610.1500 0.5200 ;
    END
  END mem_in_core0[35]
  PIN mem_in_core0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 614.0500 0.0000 614.1500 0.5200 ;
    END
  END mem_in_core0[34]
  PIN mem_in_core0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 618.0500 0.0000 618.1500 0.5200 ;
    END
  END mem_in_core0[33]
  PIN mem_in_core0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 622.0500 0.0000 622.1500 0.5200 ;
    END
  END mem_in_core0[32]
  PIN mem_in_core0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 626.0500 0.0000 626.1500 0.5200 ;
    END
  END mem_in_core0[31]
  PIN mem_in_core0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 630.0500 0.0000 630.1500 0.5200 ;
    END
  END mem_in_core0[30]
  PIN mem_in_core0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 634.0500 0.0000 634.1500 0.5200 ;
    END
  END mem_in_core0[29]
  PIN mem_in_core0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 638.0500 0.0000 638.1500 0.5200 ;
    END
  END mem_in_core0[28]
  PIN mem_in_core0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 642.0500 0.0000 642.1500 0.5200 ;
    END
  END mem_in_core0[27]
  PIN mem_in_core0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 646.0500 0.0000 646.1500 0.5200 ;
    END
  END mem_in_core0[26]
  PIN mem_in_core0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 650.0500 0.0000 650.1500 0.5200 ;
    END
  END mem_in_core0[25]
  PIN mem_in_core0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 654.0500 0.0000 654.1500 0.5200 ;
    END
  END mem_in_core0[24]
  PIN mem_in_core0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 658.0500 0.0000 658.1500 0.5200 ;
    END
  END mem_in_core0[23]
  PIN mem_in_core0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 662.0500 0.0000 662.1500 0.5200 ;
    END
  END mem_in_core0[22]
  PIN mem_in_core0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 666.0500 0.0000 666.1500 0.5200 ;
    END
  END mem_in_core0[21]
  PIN mem_in_core0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 670.0500 0.0000 670.1500 0.5200 ;
    END
  END mem_in_core0[20]
  PIN mem_in_core0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 674.0500 0.0000 674.1500 0.5200 ;
    END
  END mem_in_core0[19]
  PIN mem_in_core0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 678.0500 0.0000 678.1500 0.5200 ;
    END
  END mem_in_core0[18]
  PIN mem_in_core0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 682.0500 0.0000 682.1500 0.5200 ;
    END
  END mem_in_core0[17]
  PIN mem_in_core0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 686.0500 0.0000 686.1500 0.5200 ;
    END
  END mem_in_core0[16]
  PIN mem_in_core0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 690.0500 0.0000 690.1500 0.5200 ;
    END
  END mem_in_core0[15]
  PIN mem_in_core0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 694.0500 0.0000 694.1500 0.5200 ;
    END
  END mem_in_core0[14]
  PIN mem_in_core0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 698.0500 0.0000 698.1500 0.5200 ;
    END
  END mem_in_core0[13]
  PIN mem_in_core0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 702.0500 0.0000 702.1500 0.5200 ;
    END
  END mem_in_core0[12]
  PIN mem_in_core0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 706.0500 0.0000 706.1500 0.5200 ;
    END
  END mem_in_core0[11]
  PIN mem_in_core0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 710.0500 0.0000 710.1500 0.5200 ;
    END
  END mem_in_core0[10]
  PIN mem_in_core0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 714.0500 0.0000 714.1500 0.5200 ;
    END
  END mem_in_core0[9]
  PIN mem_in_core0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 718.0500 0.0000 718.1500 0.5200 ;
    END
  END mem_in_core0[8]
  PIN mem_in_core0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 722.0500 0.0000 722.1500 0.5200 ;
    END
  END mem_in_core0[7]
  PIN mem_in_core0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 726.0500 0.0000 726.1500 0.5200 ;
    END
  END mem_in_core0[6]
  PIN mem_in_core0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 730.0500 0.0000 730.1500 0.5200 ;
    END
  END mem_in_core0[5]
  PIN mem_in_core0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 734.0500 0.0000 734.1500 0.5200 ;
    END
  END mem_in_core0[4]
  PIN mem_in_core0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 738.0500 0.0000 738.1500 0.5200 ;
    END
  END mem_in_core0[3]
  PIN mem_in_core0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 742.0500 0.0000 742.1500 0.5200 ;
    END
  END mem_in_core0[2]
  PIN mem_in_core0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 746.0500 0.0000 746.1500 0.5200 ;
    END
  END mem_in_core0[1]
  PIN mem_in_core0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 750.0500 0.0000 750.1500 0.5200 ;
    END
  END mem_in_core0[0]
  PIN mem_in_core1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 754.0500 0.0000 754.1500 0.5200 ;
    END
  END mem_in_core1[63]
  PIN mem_in_core1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 758.0500 0.0000 758.1500 0.5200 ;
    END
  END mem_in_core1[62]
  PIN mem_in_core1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 762.0500 0.0000 762.1500 0.5200 ;
    END
  END mem_in_core1[61]
  PIN mem_in_core1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 766.0500 0.0000 766.1500 0.5200 ;
    END
  END mem_in_core1[60]
  PIN mem_in_core1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 770.0500 0.0000 770.1500 0.5200 ;
    END
  END mem_in_core1[59]
  PIN mem_in_core1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 774.0500 0.0000 774.1500 0.5200 ;
    END
  END mem_in_core1[58]
  PIN mem_in_core1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 778.0500 0.0000 778.1500 0.5200 ;
    END
  END mem_in_core1[57]
  PIN mem_in_core1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 782.0500 0.0000 782.1500 0.5200 ;
    END
  END mem_in_core1[56]
  PIN mem_in_core1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 786.0500 0.0000 786.1500 0.5200 ;
    END
  END mem_in_core1[55]
  PIN mem_in_core1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 790.0500 0.0000 790.1500 0.5200 ;
    END
  END mem_in_core1[54]
  PIN mem_in_core1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 794.0500 0.0000 794.1500 0.5200 ;
    END
  END mem_in_core1[53]
  PIN mem_in_core1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 798.0500 0.0000 798.1500 0.5200 ;
    END
  END mem_in_core1[52]
  PIN mem_in_core1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 802.0500 0.0000 802.1500 0.5200 ;
    END
  END mem_in_core1[51]
  PIN mem_in_core1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 806.0500 0.0000 806.1500 0.5200 ;
    END
  END mem_in_core1[50]
  PIN mem_in_core1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 810.0500 0.0000 810.1500 0.5200 ;
    END
  END mem_in_core1[49]
  PIN mem_in_core1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 814.0500 0.0000 814.1500 0.5200 ;
    END
  END mem_in_core1[48]
  PIN mem_in_core1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 818.0500 0.0000 818.1500 0.5200 ;
    END
  END mem_in_core1[47]
  PIN mem_in_core1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 822.0500 0.0000 822.1500 0.5200 ;
    END
  END mem_in_core1[46]
  PIN mem_in_core1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 826.0500 0.0000 826.1500 0.5200 ;
    END
  END mem_in_core1[45]
  PIN mem_in_core1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 830.0500 0.0000 830.1500 0.5200 ;
    END
  END mem_in_core1[44]
  PIN mem_in_core1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 834.0500 0.0000 834.1500 0.5200 ;
    END
  END mem_in_core1[43]
  PIN mem_in_core1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 838.0500 0.0000 838.1500 0.5200 ;
    END
  END mem_in_core1[42]
  PIN mem_in_core1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 842.0500 0.0000 842.1500 0.5200 ;
    END
  END mem_in_core1[41]
  PIN mem_in_core1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 846.0500 0.0000 846.1500 0.5200 ;
    END
  END mem_in_core1[40]
  PIN mem_in_core1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 850.0500 0.0000 850.1500 0.5200 ;
    END
  END mem_in_core1[39]
  PIN mem_in_core1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 854.0500 0.0000 854.1500 0.5200 ;
    END
  END mem_in_core1[38]
  PIN mem_in_core1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 858.0500 0.0000 858.1500 0.5200 ;
    END
  END mem_in_core1[37]
  PIN mem_in_core1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 862.0500 0.0000 862.1500 0.5200 ;
    END
  END mem_in_core1[36]
  PIN mem_in_core1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 866.0500 0.0000 866.1500 0.5200 ;
    END
  END mem_in_core1[35]
  PIN mem_in_core1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 870.0500 0.0000 870.1500 0.5200 ;
    END
  END mem_in_core1[34]
  PIN mem_in_core1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 874.0500 0.0000 874.1500 0.5200 ;
    END
  END mem_in_core1[33]
  PIN mem_in_core1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 878.0500 0.0000 878.1500 0.5200 ;
    END
  END mem_in_core1[32]
  PIN mem_in_core1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 882.0500 0.0000 882.1500 0.5200 ;
    END
  END mem_in_core1[31]
  PIN mem_in_core1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 886.0500 0.0000 886.1500 0.5200 ;
    END
  END mem_in_core1[30]
  PIN mem_in_core1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 890.0500 0.0000 890.1500 0.5200 ;
    END
  END mem_in_core1[29]
  PIN mem_in_core1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 894.0500 0.0000 894.1500 0.5200 ;
    END
  END mem_in_core1[28]
  PIN mem_in_core1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 898.0500 0.0000 898.1500 0.5200 ;
    END
  END mem_in_core1[27]
  PIN mem_in_core1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 902.0500 0.0000 902.1500 0.5200 ;
    END
  END mem_in_core1[26]
  PIN mem_in_core1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 906.0500 0.0000 906.1500 0.5200 ;
    END
  END mem_in_core1[25]
  PIN mem_in_core1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 910.0500 0.0000 910.1500 0.5200 ;
    END
  END mem_in_core1[24]
  PIN mem_in_core1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 914.0500 0.0000 914.1500 0.5200 ;
    END
  END mem_in_core1[23]
  PIN mem_in_core1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 918.0500 0.0000 918.1500 0.5200 ;
    END
  END mem_in_core1[22]
  PIN mem_in_core1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 922.0500 0.0000 922.1500 0.5200 ;
    END
  END mem_in_core1[21]
  PIN mem_in_core1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 926.0500 0.0000 926.1500 0.5200 ;
    END
  END mem_in_core1[20]
  PIN mem_in_core1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 930.0500 0.0000 930.1500 0.5200 ;
    END
  END mem_in_core1[19]
  PIN mem_in_core1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 934.0500 0.0000 934.1500 0.5200 ;
    END
  END mem_in_core1[18]
  PIN mem_in_core1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 938.0500 0.0000 938.1500 0.5200 ;
    END
  END mem_in_core1[17]
  PIN mem_in_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 942.0500 0.0000 942.1500 0.5200 ;
    END
  END mem_in_core1[16]
  PIN mem_in_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 946.0500 0.0000 946.1500 0.5200 ;
    END
  END mem_in_core1[15]
  PIN mem_in_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 950.0500 0.0000 950.1500 0.5200 ;
    END
  END mem_in_core1[14]
  PIN mem_in_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 954.0500 0.0000 954.1500 0.5200 ;
    END
  END mem_in_core1[13]
  PIN mem_in_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 958.0500 0.0000 958.1500 0.5200 ;
    END
  END mem_in_core1[12]
  PIN mem_in_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 962.0500 0.0000 962.1500 0.5200 ;
    END
  END mem_in_core1[11]
  PIN mem_in_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 966.0500 0.0000 966.1500 0.5200 ;
    END
  END mem_in_core1[10]
  PIN mem_in_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 970.0500 0.0000 970.1500 0.5200 ;
    END
  END mem_in_core1[9]
  PIN mem_in_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 974.0500 0.0000 974.1500 0.5200 ;
    END
  END mem_in_core1[8]
  PIN mem_in_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 978.0500 0.0000 978.1500 0.5200 ;
    END
  END mem_in_core1[7]
  PIN mem_in_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 982.0500 0.0000 982.1500 0.5200 ;
    END
  END mem_in_core1[6]
  PIN mem_in_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 986.0500 0.0000 986.1500 0.5200 ;
    END
  END mem_in_core1[5]
  PIN mem_in_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 990.0500 0.0000 990.1500 0.5200 ;
    END
  END mem_in_core1[4]
  PIN mem_in_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 994.0500 0.0000 994.1500 0.5200 ;
    END
  END mem_in_core1[3]
  PIN mem_in_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 998.0500 0.0000 998.1500 0.5200 ;
    END
  END mem_in_core1[2]
  PIN mem_in_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1002.0500 0.0000 1002.1500 0.5200 ;
    END
  END mem_in_core1[1]
  PIN mem_in_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1006.0500 0.0000 1006.1500 0.5200 ;
    END
  END mem_in_core1[0]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 422.0500 0.0000 422.1500 0.5200 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 426.0500 0.0000 426.1500 0.5200 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 430.0500 0.0000 430.1500 0.5200 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 434.0500 0.0000 434.1500 0.5200 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 438.0500 0.0000 438.1500 0.5200 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 442.0500 0.0000 442.1500 0.5200 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 446.0500 0.0000 446.1500 0.5200 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 450.0500 0.0000 450.1500 0.5200 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 454.0500 0.0000 454.1500 0.5200 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 458.0500 0.0000 458.1500 0.5200 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 462.0500 0.0000 462.1500 0.5200 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 466.0500 0.0000 466.1500 0.5200 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 470.0500 0.0000 470.1500 0.5200 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 474.0500 0.0000 474.1500 0.5200 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 478.0500 0.0000 478.1500 0.5200 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 482.0500 0.0000 482.1500 0.5200 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 486.0500 0.0000 486.1500 0.5200 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 490.0500 0.0000 490.1500 0.5200 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 494.0500 0.0000 494.1500 0.5200 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 414.0500 0.0000 414.1500 0.5200 ;
    END
  END reset
  PIN out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1347.8500 2819.4800 1347.9500 2820.0000 ;
    END
  END out[319]
  PIN out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1343.8500 2819.4800 1343.9500 2820.0000 ;
    END
  END out[318]
  PIN out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1339.8500 2819.4800 1339.9500 2820.0000 ;
    END
  END out[317]
  PIN out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1335.8500 2819.4800 1335.9500 2820.0000 ;
    END
  END out[316]
  PIN out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1331.8500 2819.4800 1331.9500 2820.0000 ;
    END
  END out[315]
  PIN out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1327.8500 2819.4800 1327.9500 2820.0000 ;
    END
  END out[314]
  PIN out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1323.8500 2819.4800 1323.9500 2820.0000 ;
    END
  END out[313]
  PIN out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1319.8500 2819.4800 1319.9500 2820.0000 ;
    END
  END out[312]
  PIN out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1315.8500 2819.4800 1315.9500 2820.0000 ;
    END
  END out[311]
  PIN out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1311.8500 2819.4800 1311.9500 2820.0000 ;
    END
  END out[310]
  PIN out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1307.8500 2819.4800 1307.9500 2820.0000 ;
    END
  END out[309]
  PIN out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1303.8500 2819.4800 1303.9500 2820.0000 ;
    END
  END out[308]
  PIN out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1299.8500 2819.4800 1299.9500 2820.0000 ;
    END
  END out[307]
  PIN out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1295.8500 2819.4800 1295.9500 2820.0000 ;
    END
  END out[306]
  PIN out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1291.8500 2819.4800 1291.9500 2820.0000 ;
    END
  END out[305]
  PIN out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1287.8500 2819.4800 1287.9500 2820.0000 ;
    END
  END out[304]
  PIN out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1283.8500 2819.4800 1283.9500 2820.0000 ;
    END
  END out[303]
  PIN out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1279.8500 2819.4800 1279.9500 2820.0000 ;
    END
  END out[302]
  PIN out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1275.8500 2819.4800 1275.9500 2820.0000 ;
    END
  END out[301]
  PIN out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1271.8500 2819.4800 1271.9500 2820.0000 ;
    END
  END out[300]
  PIN out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1267.8500 2819.4800 1267.9500 2820.0000 ;
    END
  END out[299]
  PIN out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1263.8500 2819.4800 1263.9500 2820.0000 ;
    END
  END out[298]
  PIN out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1259.8500 2819.4800 1259.9500 2820.0000 ;
    END
  END out[297]
  PIN out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1255.8500 2819.4800 1255.9500 2820.0000 ;
    END
  END out[296]
  PIN out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1251.8500 2819.4800 1251.9500 2820.0000 ;
    END
  END out[295]
  PIN out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1247.8500 2819.4800 1247.9500 2820.0000 ;
    END
  END out[294]
  PIN out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1243.8500 2819.4800 1243.9500 2820.0000 ;
    END
  END out[293]
  PIN out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1239.8500 2819.4800 1239.9500 2820.0000 ;
    END
  END out[292]
  PIN out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1235.8500 2819.4800 1235.9500 2820.0000 ;
    END
  END out[291]
  PIN out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1231.8500 2819.4800 1231.9500 2820.0000 ;
    END
  END out[290]
  PIN out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1227.8500 2819.4800 1227.9500 2820.0000 ;
    END
  END out[289]
  PIN out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1223.8500 2819.4800 1223.9500 2820.0000 ;
    END
  END out[288]
  PIN out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1219.8500 2819.4800 1219.9500 2820.0000 ;
    END
  END out[287]
  PIN out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1215.8500 2819.4800 1215.9500 2820.0000 ;
    END
  END out[286]
  PIN out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1211.8500 2819.4800 1211.9500 2820.0000 ;
    END
  END out[285]
  PIN out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1207.8500 2819.4800 1207.9500 2820.0000 ;
    END
  END out[284]
  PIN out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1203.8500 2819.4800 1203.9500 2820.0000 ;
    END
  END out[283]
  PIN out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1199.8500 2819.4800 1199.9500 2820.0000 ;
    END
  END out[282]
  PIN out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1195.8500 2819.4800 1195.9500 2820.0000 ;
    END
  END out[281]
  PIN out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1191.8500 2819.4800 1191.9500 2820.0000 ;
    END
  END out[280]
  PIN out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1187.8500 2819.4800 1187.9500 2820.0000 ;
    END
  END out[279]
  PIN out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1183.8500 2819.4800 1183.9500 2820.0000 ;
    END
  END out[278]
  PIN out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1179.8500 2819.4800 1179.9500 2820.0000 ;
    END
  END out[277]
  PIN out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1175.8500 2819.4800 1175.9500 2820.0000 ;
    END
  END out[276]
  PIN out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1171.8500 2819.4800 1171.9500 2820.0000 ;
    END
  END out[275]
  PIN out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1167.8500 2819.4800 1167.9500 2820.0000 ;
    END
  END out[274]
  PIN out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1163.8500 2819.4800 1163.9500 2820.0000 ;
    END
  END out[273]
  PIN out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1159.8500 2819.4800 1159.9500 2820.0000 ;
    END
  END out[272]
  PIN out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1155.8500 2819.4800 1155.9500 2820.0000 ;
    END
  END out[271]
  PIN out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1151.8500 2819.4800 1151.9500 2820.0000 ;
    END
  END out[270]
  PIN out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1147.8500 2819.4800 1147.9500 2820.0000 ;
    END
  END out[269]
  PIN out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1143.8500 2819.4800 1143.9500 2820.0000 ;
    END
  END out[268]
  PIN out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1139.8500 2819.4800 1139.9500 2820.0000 ;
    END
  END out[267]
  PIN out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1135.8500 2819.4800 1135.9500 2820.0000 ;
    END
  END out[266]
  PIN out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1131.8500 2819.4800 1131.9500 2820.0000 ;
    END
  END out[265]
  PIN out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1127.8500 2819.4800 1127.9500 2820.0000 ;
    END
  END out[264]
  PIN out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1123.8500 2819.4800 1123.9500 2820.0000 ;
    END
  END out[263]
  PIN out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1119.8500 2819.4800 1119.9500 2820.0000 ;
    END
  END out[262]
  PIN out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1115.8500 2819.4800 1115.9500 2820.0000 ;
    END
  END out[261]
  PIN out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1111.8500 2819.4800 1111.9500 2820.0000 ;
    END
  END out[260]
  PIN out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1107.8500 2819.4800 1107.9500 2820.0000 ;
    END
  END out[259]
  PIN out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1103.8500 2819.4800 1103.9500 2820.0000 ;
    END
  END out[258]
  PIN out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1099.8500 2819.4800 1099.9500 2820.0000 ;
    END
  END out[257]
  PIN out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1095.8500 2819.4800 1095.9500 2820.0000 ;
    END
  END out[256]
  PIN out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1091.8500 2819.4800 1091.9500 2820.0000 ;
    END
  END out[255]
  PIN out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1087.8500 2819.4800 1087.9500 2820.0000 ;
    END
  END out[254]
  PIN out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1083.8500 2819.4800 1083.9500 2820.0000 ;
    END
  END out[253]
  PIN out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1079.8500 2819.4800 1079.9500 2820.0000 ;
    END
  END out[252]
  PIN out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1075.8500 2819.4800 1075.9500 2820.0000 ;
    END
  END out[251]
  PIN out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1071.8500 2819.4800 1071.9500 2820.0000 ;
    END
  END out[250]
  PIN out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1067.8500 2819.4800 1067.9500 2820.0000 ;
    END
  END out[249]
  PIN out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1063.8500 2819.4800 1063.9500 2820.0000 ;
    END
  END out[248]
  PIN out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1059.8500 2819.4800 1059.9500 2820.0000 ;
    END
  END out[247]
  PIN out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1055.8500 2819.4800 1055.9500 2820.0000 ;
    END
  END out[246]
  PIN out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1051.8500 2819.4800 1051.9500 2820.0000 ;
    END
  END out[245]
  PIN out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1047.8500 2819.4800 1047.9500 2820.0000 ;
    END
  END out[244]
  PIN out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1043.8500 2819.4800 1043.9500 2820.0000 ;
    END
  END out[243]
  PIN out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1039.8500 2819.4800 1039.9500 2820.0000 ;
    END
  END out[242]
  PIN out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1035.8500 2819.4800 1035.9500 2820.0000 ;
    END
  END out[241]
  PIN out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1031.8500 2819.4800 1031.9500 2820.0000 ;
    END
  END out[240]
  PIN out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1027.8500 2819.4800 1027.9500 2820.0000 ;
    END
  END out[239]
  PIN out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1023.8500 2819.4800 1023.9500 2820.0000 ;
    END
  END out[238]
  PIN out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1019.8500 2819.4800 1019.9500 2820.0000 ;
    END
  END out[237]
  PIN out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1015.8500 2819.4800 1015.9500 2820.0000 ;
    END
  END out[236]
  PIN out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1011.8500 2819.4800 1011.9500 2820.0000 ;
    END
  END out[235]
  PIN out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1007.8500 2819.4800 1007.9500 2820.0000 ;
    END
  END out[234]
  PIN out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1003.8500 2819.4800 1003.9500 2820.0000 ;
    END
  END out[233]
  PIN out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 999.8500 2819.4800 999.9500 2820.0000 ;
    END
  END out[232]
  PIN out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 995.8500 2819.4800 995.9500 2820.0000 ;
    END
  END out[231]
  PIN out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 991.8500 2819.4800 991.9500 2820.0000 ;
    END
  END out[230]
  PIN out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 987.8500 2819.4800 987.9500 2820.0000 ;
    END
  END out[229]
  PIN out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 983.8500 2819.4800 983.9500 2820.0000 ;
    END
  END out[228]
  PIN out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 979.8500 2819.4800 979.9500 2820.0000 ;
    END
  END out[227]
  PIN out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 975.8500 2819.4800 975.9500 2820.0000 ;
    END
  END out[226]
  PIN out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 971.8500 2819.4800 971.9500 2820.0000 ;
    END
  END out[225]
  PIN out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 967.8500 2819.4800 967.9500 2820.0000 ;
    END
  END out[224]
  PIN out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 963.8500 2819.4800 963.9500 2820.0000 ;
    END
  END out[223]
  PIN out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 959.8500 2819.4800 959.9500 2820.0000 ;
    END
  END out[222]
  PIN out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 955.8500 2819.4800 955.9500 2820.0000 ;
    END
  END out[221]
  PIN out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 951.8500 2819.4800 951.9500 2820.0000 ;
    END
  END out[220]
  PIN out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 947.8500 2819.4800 947.9500 2820.0000 ;
    END
  END out[219]
  PIN out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 943.8500 2819.4800 943.9500 2820.0000 ;
    END
  END out[218]
  PIN out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 939.8500 2819.4800 939.9500 2820.0000 ;
    END
  END out[217]
  PIN out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 935.8500 2819.4800 935.9500 2820.0000 ;
    END
  END out[216]
  PIN out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 931.8500 2819.4800 931.9500 2820.0000 ;
    END
  END out[215]
  PIN out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 927.8500 2819.4800 927.9500 2820.0000 ;
    END
  END out[214]
  PIN out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 923.8500 2819.4800 923.9500 2820.0000 ;
    END
  END out[213]
  PIN out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 919.8500 2819.4800 919.9500 2820.0000 ;
    END
  END out[212]
  PIN out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 915.8500 2819.4800 915.9500 2820.0000 ;
    END
  END out[211]
  PIN out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 911.8500 2819.4800 911.9500 2820.0000 ;
    END
  END out[210]
  PIN out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 907.8500 2819.4800 907.9500 2820.0000 ;
    END
  END out[209]
  PIN out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 903.8500 2819.4800 903.9500 2820.0000 ;
    END
  END out[208]
  PIN out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 899.8500 2819.4800 899.9500 2820.0000 ;
    END
  END out[207]
  PIN out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 895.8500 2819.4800 895.9500 2820.0000 ;
    END
  END out[206]
  PIN out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 891.8500 2819.4800 891.9500 2820.0000 ;
    END
  END out[205]
  PIN out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 887.8500 2819.4800 887.9500 2820.0000 ;
    END
  END out[204]
  PIN out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 883.8500 2819.4800 883.9500 2820.0000 ;
    END
  END out[203]
  PIN out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 879.8500 2819.4800 879.9500 2820.0000 ;
    END
  END out[202]
  PIN out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 875.8500 2819.4800 875.9500 2820.0000 ;
    END
  END out[201]
  PIN out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 871.8500 2819.4800 871.9500 2820.0000 ;
    END
  END out[200]
  PIN out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 867.8500 2819.4800 867.9500 2820.0000 ;
    END
  END out[199]
  PIN out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 863.8500 2819.4800 863.9500 2820.0000 ;
    END
  END out[198]
  PIN out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 859.8500 2819.4800 859.9500 2820.0000 ;
    END
  END out[197]
  PIN out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 855.8500 2819.4800 855.9500 2820.0000 ;
    END
  END out[196]
  PIN out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 851.8500 2819.4800 851.9500 2820.0000 ;
    END
  END out[195]
  PIN out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 847.8500 2819.4800 847.9500 2820.0000 ;
    END
  END out[194]
  PIN out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 843.8500 2819.4800 843.9500 2820.0000 ;
    END
  END out[193]
  PIN out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 839.8500 2819.4800 839.9500 2820.0000 ;
    END
  END out[192]
  PIN out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 835.8500 2819.4800 835.9500 2820.0000 ;
    END
  END out[191]
  PIN out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 831.8500 2819.4800 831.9500 2820.0000 ;
    END
  END out[190]
  PIN out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 827.8500 2819.4800 827.9500 2820.0000 ;
    END
  END out[189]
  PIN out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 823.8500 2819.4800 823.9500 2820.0000 ;
    END
  END out[188]
  PIN out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 819.8500 2819.4800 819.9500 2820.0000 ;
    END
  END out[187]
  PIN out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 815.8500 2819.4800 815.9500 2820.0000 ;
    END
  END out[186]
  PIN out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 811.8500 2819.4800 811.9500 2820.0000 ;
    END
  END out[185]
  PIN out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 807.8500 2819.4800 807.9500 2820.0000 ;
    END
  END out[184]
  PIN out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 803.8500 2819.4800 803.9500 2820.0000 ;
    END
  END out[183]
  PIN out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 799.8500 2819.4800 799.9500 2820.0000 ;
    END
  END out[182]
  PIN out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 795.8500 2819.4800 795.9500 2820.0000 ;
    END
  END out[181]
  PIN out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 791.8500 2819.4800 791.9500 2820.0000 ;
    END
  END out[180]
  PIN out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 787.8500 2819.4800 787.9500 2820.0000 ;
    END
  END out[179]
  PIN out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 783.8500 2819.4800 783.9500 2820.0000 ;
    END
  END out[178]
  PIN out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 779.8500 2819.4800 779.9500 2820.0000 ;
    END
  END out[177]
  PIN out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 775.8500 2819.4800 775.9500 2820.0000 ;
    END
  END out[176]
  PIN out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 771.8500 2819.4800 771.9500 2820.0000 ;
    END
  END out[175]
  PIN out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 767.8500 2819.4800 767.9500 2820.0000 ;
    END
  END out[174]
  PIN out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 763.8500 2819.4800 763.9500 2820.0000 ;
    END
  END out[173]
  PIN out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 759.8500 2819.4800 759.9500 2820.0000 ;
    END
  END out[172]
  PIN out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 755.8500 2819.4800 755.9500 2820.0000 ;
    END
  END out[171]
  PIN out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 751.8500 2819.4800 751.9500 2820.0000 ;
    END
  END out[170]
  PIN out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 747.8500 2819.4800 747.9500 2820.0000 ;
    END
  END out[169]
  PIN out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 743.8500 2819.4800 743.9500 2820.0000 ;
    END
  END out[168]
  PIN out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 739.8500 2819.4800 739.9500 2820.0000 ;
    END
  END out[167]
  PIN out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 735.8500 2819.4800 735.9500 2820.0000 ;
    END
  END out[166]
  PIN out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 731.8500 2819.4800 731.9500 2820.0000 ;
    END
  END out[165]
  PIN out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 727.8500 2819.4800 727.9500 2820.0000 ;
    END
  END out[164]
  PIN out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 723.8500 2819.4800 723.9500 2820.0000 ;
    END
  END out[163]
  PIN out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 719.8500 2819.4800 719.9500 2820.0000 ;
    END
  END out[162]
  PIN out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 715.8500 2819.4800 715.9500 2820.0000 ;
    END
  END out[161]
  PIN out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 711.8500 2819.4800 711.9500 2820.0000 ;
    END
  END out[160]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 707.8500 2819.4800 707.9500 2820.0000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 703.8500 2819.4800 703.9500 2820.0000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 699.8500 2819.4800 699.9500 2820.0000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 695.8500 2819.4800 695.9500 2820.0000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 691.8500 2819.4800 691.9500 2820.0000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 687.8500 2819.4800 687.9500 2820.0000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 683.8500 2819.4800 683.9500 2820.0000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 679.8500 2819.4800 679.9500 2820.0000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 675.8500 2819.4800 675.9500 2820.0000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 671.8500 2819.4800 671.9500 2820.0000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 667.8500 2819.4800 667.9500 2820.0000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 663.8500 2819.4800 663.9500 2820.0000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 659.8500 2819.4800 659.9500 2820.0000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 655.8500 2819.4800 655.9500 2820.0000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 651.8500 2819.4800 651.9500 2820.0000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 647.8500 2819.4800 647.9500 2820.0000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 643.8500 2819.4800 643.9500 2820.0000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 639.8500 2819.4800 639.9500 2820.0000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 635.8500 2819.4800 635.9500 2820.0000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 631.8500 2819.4800 631.9500 2820.0000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 627.8500 2819.4800 627.9500 2820.0000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 623.8500 2819.4800 623.9500 2820.0000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 619.8500 2819.4800 619.9500 2820.0000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 615.8500 2819.4800 615.9500 2820.0000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 611.8500 2819.4800 611.9500 2820.0000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 607.8500 2819.4800 607.9500 2820.0000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 603.8500 2819.4800 603.9500 2820.0000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 599.8500 2819.4800 599.9500 2820.0000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 595.8500 2819.4800 595.9500 2820.0000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 591.8500 2819.4800 591.9500 2820.0000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 587.8500 2819.4800 587.9500 2820.0000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 583.8500 2819.4800 583.9500 2820.0000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 579.8500 2819.4800 579.9500 2820.0000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 575.8500 2819.4800 575.9500 2820.0000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 571.8500 2819.4800 571.9500 2820.0000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 567.8500 2819.4800 567.9500 2820.0000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 563.8500 2819.4800 563.9500 2820.0000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 559.8500 2819.4800 559.9500 2820.0000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 555.8500 2819.4800 555.9500 2820.0000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 551.8500 2819.4800 551.9500 2820.0000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 547.8500 2819.4800 547.9500 2820.0000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 543.8500 2819.4800 543.9500 2820.0000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 539.8500 2819.4800 539.9500 2820.0000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 535.8500 2819.4800 535.9500 2820.0000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 531.8500 2819.4800 531.9500 2820.0000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 527.8500 2819.4800 527.9500 2820.0000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 523.8500 2819.4800 523.9500 2820.0000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 519.8500 2819.4800 519.9500 2820.0000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 515.8500 2819.4800 515.9500 2820.0000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 511.8500 2819.4800 511.9500 2820.0000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 507.8500 2819.4800 507.9500 2820.0000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 503.8500 2819.4800 503.9500 2820.0000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 499.8500 2819.4800 499.9500 2820.0000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 495.8500 2819.4800 495.9500 2820.0000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 491.8500 2819.4800 491.9500 2820.0000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 487.8500 2819.4800 487.9500 2820.0000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 483.8500 2819.4800 483.9500 2820.0000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 479.8500 2819.4800 479.9500 2820.0000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 475.8500 2819.4800 475.9500 2820.0000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 471.8500 2819.4800 471.9500 2820.0000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 467.8500 2819.4800 467.9500 2820.0000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 463.8500 2819.4800 463.9500 2820.0000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 459.8500 2819.4800 459.9500 2820.0000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 455.8500 2819.4800 455.9500 2820.0000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 451.8500 2819.4800 451.9500 2820.0000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 447.8500 2819.4800 447.9500 2820.0000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 443.8500 2819.4800 443.9500 2820.0000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 439.8500 2819.4800 439.9500 2820.0000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 435.8500 2819.4800 435.9500 2820.0000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 431.8500 2819.4800 431.9500 2820.0000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 427.8500 2819.4800 427.9500 2820.0000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 423.8500 2819.4800 423.9500 2820.0000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 419.8500 2819.4800 419.9500 2820.0000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 415.8500 2819.4800 415.9500 2820.0000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 411.8500 2819.4800 411.9500 2820.0000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 407.8500 2819.4800 407.9500 2820.0000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 403.8500 2819.4800 403.9500 2820.0000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 399.8500 2819.4800 399.9500 2820.0000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 395.8500 2819.4800 395.9500 2820.0000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 391.8500 2819.4800 391.9500 2820.0000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 387.8500 2819.4800 387.9500 2820.0000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 383.8500 2819.4800 383.9500 2820.0000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 379.8500 2819.4800 379.9500 2820.0000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 375.8500 2819.4800 375.9500 2820.0000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 371.8500 2819.4800 371.9500 2820.0000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 367.8500 2819.4800 367.9500 2820.0000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 363.8500 2819.4800 363.9500 2820.0000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 359.8500 2819.4800 359.9500 2820.0000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 355.8500 2819.4800 355.9500 2820.0000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 351.8500 2819.4800 351.9500 2820.0000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 347.8500 2819.4800 347.9500 2820.0000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 343.8500 2819.4800 343.9500 2820.0000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 339.8500 2819.4800 339.9500 2820.0000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 335.8500 2819.4800 335.9500 2820.0000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 331.8500 2819.4800 331.9500 2820.0000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 327.8500 2819.4800 327.9500 2820.0000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 323.8500 2819.4800 323.9500 2820.0000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 319.8500 2819.4800 319.9500 2820.0000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 315.8500 2819.4800 315.9500 2820.0000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 311.8500 2819.4800 311.9500 2820.0000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 307.8500 2819.4800 307.9500 2820.0000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 303.8500 2819.4800 303.9500 2820.0000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 299.8500 2819.4800 299.9500 2820.0000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 295.8500 2819.4800 295.9500 2820.0000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 291.8500 2819.4800 291.9500 2820.0000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 287.8500 2819.4800 287.9500 2820.0000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 283.8500 2819.4800 283.9500 2820.0000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 279.8500 2819.4800 279.9500 2820.0000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 275.8500 2819.4800 275.9500 2820.0000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 271.8500 2819.4800 271.9500 2820.0000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 267.8500 2819.4800 267.9500 2820.0000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 263.8500 2819.4800 263.9500 2820.0000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 259.8500 2819.4800 259.9500 2820.0000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 255.8500 2819.4800 255.9500 2820.0000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 251.8500 2819.4800 251.9500 2820.0000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 247.8500 2819.4800 247.9500 2820.0000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 243.8500 2819.4800 243.9500 2820.0000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 239.8500 2819.4800 239.9500 2820.0000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 235.8500 2819.4800 235.9500 2820.0000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 231.8500 2819.4800 231.9500 2820.0000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 227.8500 2819.4800 227.9500 2820.0000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 223.8500 2819.4800 223.9500 2820.0000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 219.8500 2819.4800 219.9500 2820.0000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 215.8500 2819.4800 215.9500 2820.0000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 211.8500 2819.4800 211.9500 2820.0000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 207.8500 2819.4800 207.9500 2820.0000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 203.8500 2819.4800 203.9500 2820.0000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 199.8500 2819.4800 199.9500 2820.0000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 195.8500 2819.4800 195.9500 2820.0000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 191.8500 2819.4800 191.9500 2820.0000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 187.8500 2819.4800 187.9500 2820.0000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 183.8500 2819.4800 183.9500 2820.0000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 179.8500 2819.4800 179.9500 2820.0000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 175.8500 2819.4800 175.9500 2820.0000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 171.8500 2819.4800 171.9500 2820.0000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 167.8500 2819.4800 167.9500 2820.0000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 163.8500 2819.4800 163.9500 2820.0000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 159.8500 2819.4800 159.9500 2820.0000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 155.8500 2819.4800 155.9500 2820.0000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 151.8500 2819.4800 151.9500 2820.0000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 147.8500 2819.4800 147.9500 2820.0000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 143.8500 2819.4800 143.9500 2820.0000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 139.8500 2819.4800 139.9500 2820.0000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 135.8500 2819.4800 135.9500 2820.0000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 131.8500 2819.4800 131.9500 2820.0000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 127.8500 2819.4800 127.9500 2820.0000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 123.8500 2819.4800 123.9500 2820.0000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 119.8500 2819.4800 119.9500 2820.0000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 115.8500 2819.4800 115.9500 2820.0000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 111.8500 2819.4800 111.9500 2820.0000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 107.8500 2819.4800 107.9500 2820.0000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 103.8500 2819.4800 103.9500 2820.0000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 99.8500 2819.4800 99.9500 2820.0000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 95.8500 2819.4800 95.9500 2820.0000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 91.8500 2819.4800 91.9500 2820.0000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 87.8500 2819.4800 87.9500 2820.0000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 83.8500 2819.4800 83.9500 2820.0000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 79.8500 2819.4800 79.9500 2820.0000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 75.8500 2819.4800 75.9500 2820.0000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 71.8500 2819.4800 71.9500 2820.0000 ;
    END
  END out[0]
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M4 ;
      RECT 1348.0500 2819.3800 1420.0000 2820.0000 ;
      RECT 1344.0500 2819.3800 1347.7500 2820.0000 ;
      RECT 1340.0500 2819.3800 1343.7500 2820.0000 ;
      RECT 1336.0500 2819.3800 1339.7500 2820.0000 ;
      RECT 1332.0500 2819.3800 1335.7500 2820.0000 ;
      RECT 1328.0500 2819.3800 1331.7500 2820.0000 ;
      RECT 1324.0500 2819.3800 1327.7500 2820.0000 ;
      RECT 1320.0500 2819.3800 1323.7500 2820.0000 ;
      RECT 1316.0500 2819.3800 1319.7500 2820.0000 ;
      RECT 1312.0500 2819.3800 1315.7500 2820.0000 ;
      RECT 1308.0500 2819.3800 1311.7500 2820.0000 ;
      RECT 1304.0500 2819.3800 1307.7500 2820.0000 ;
      RECT 1300.0500 2819.3800 1303.7500 2820.0000 ;
      RECT 1296.0500 2819.3800 1299.7500 2820.0000 ;
      RECT 1292.0500 2819.3800 1295.7500 2820.0000 ;
      RECT 1288.0500 2819.3800 1291.7500 2820.0000 ;
      RECT 1284.0500 2819.3800 1287.7500 2820.0000 ;
      RECT 1280.0500 2819.3800 1283.7500 2820.0000 ;
      RECT 1276.0500 2819.3800 1279.7500 2820.0000 ;
      RECT 1272.0500 2819.3800 1275.7500 2820.0000 ;
      RECT 1268.0500 2819.3800 1271.7500 2820.0000 ;
      RECT 1264.0500 2819.3800 1267.7500 2820.0000 ;
      RECT 1260.0500 2819.3800 1263.7500 2820.0000 ;
      RECT 1256.0500 2819.3800 1259.7500 2820.0000 ;
      RECT 1252.0500 2819.3800 1255.7500 2820.0000 ;
      RECT 1248.0500 2819.3800 1251.7500 2820.0000 ;
      RECT 1244.0500 2819.3800 1247.7500 2820.0000 ;
      RECT 1240.0500 2819.3800 1243.7500 2820.0000 ;
      RECT 1236.0500 2819.3800 1239.7500 2820.0000 ;
      RECT 1232.0500 2819.3800 1235.7500 2820.0000 ;
      RECT 1228.0500 2819.3800 1231.7500 2820.0000 ;
      RECT 1224.0500 2819.3800 1227.7500 2820.0000 ;
      RECT 1220.0500 2819.3800 1223.7500 2820.0000 ;
      RECT 1216.0500 2819.3800 1219.7500 2820.0000 ;
      RECT 1212.0500 2819.3800 1215.7500 2820.0000 ;
      RECT 1208.0500 2819.3800 1211.7500 2820.0000 ;
      RECT 1204.0500 2819.3800 1207.7500 2820.0000 ;
      RECT 1200.0500 2819.3800 1203.7500 2820.0000 ;
      RECT 1196.0500 2819.3800 1199.7500 2820.0000 ;
      RECT 1192.0500 2819.3800 1195.7500 2820.0000 ;
      RECT 1188.0500 2819.3800 1191.7500 2820.0000 ;
      RECT 1184.0500 2819.3800 1187.7500 2820.0000 ;
      RECT 1180.0500 2819.3800 1183.7500 2820.0000 ;
      RECT 1176.0500 2819.3800 1179.7500 2820.0000 ;
      RECT 1172.0500 2819.3800 1175.7500 2820.0000 ;
      RECT 1168.0500 2819.3800 1171.7500 2820.0000 ;
      RECT 1164.0500 2819.3800 1167.7500 2820.0000 ;
      RECT 1160.0500 2819.3800 1163.7500 2820.0000 ;
      RECT 1156.0500 2819.3800 1159.7500 2820.0000 ;
      RECT 1152.0500 2819.3800 1155.7500 2820.0000 ;
      RECT 1148.0500 2819.3800 1151.7500 2820.0000 ;
      RECT 1144.0500 2819.3800 1147.7500 2820.0000 ;
      RECT 1140.0500 2819.3800 1143.7500 2820.0000 ;
      RECT 1136.0500 2819.3800 1139.7500 2820.0000 ;
      RECT 1132.0500 2819.3800 1135.7500 2820.0000 ;
      RECT 1128.0500 2819.3800 1131.7500 2820.0000 ;
      RECT 1124.0500 2819.3800 1127.7500 2820.0000 ;
      RECT 1120.0500 2819.3800 1123.7500 2820.0000 ;
      RECT 1116.0500 2819.3800 1119.7500 2820.0000 ;
      RECT 1112.0500 2819.3800 1115.7500 2820.0000 ;
      RECT 1108.0500 2819.3800 1111.7500 2820.0000 ;
      RECT 1104.0500 2819.3800 1107.7500 2820.0000 ;
      RECT 1100.0500 2819.3800 1103.7500 2820.0000 ;
      RECT 1096.0500 2819.3800 1099.7500 2820.0000 ;
      RECT 1092.0500 2819.3800 1095.7500 2820.0000 ;
      RECT 1088.0500 2819.3800 1091.7500 2820.0000 ;
      RECT 1084.0500 2819.3800 1087.7500 2820.0000 ;
      RECT 1080.0500 2819.3800 1083.7500 2820.0000 ;
      RECT 1076.0500 2819.3800 1079.7500 2820.0000 ;
      RECT 1072.0500 2819.3800 1075.7500 2820.0000 ;
      RECT 1068.0500 2819.3800 1071.7500 2820.0000 ;
      RECT 1064.0500 2819.3800 1067.7500 2820.0000 ;
      RECT 1060.0500 2819.3800 1063.7500 2820.0000 ;
      RECT 1056.0500 2819.3800 1059.7500 2820.0000 ;
      RECT 1052.0500 2819.3800 1055.7500 2820.0000 ;
      RECT 1048.0500 2819.3800 1051.7500 2820.0000 ;
      RECT 1044.0500 2819.3800 1047.7500 2820.0000 ;
      RECT 1040.0500 2819.3800 1043.7500 2820.0000 ;
      RECT 1036.0500 2819.3800 1039.7500 2820.0000 ;
      RECT 1032.0500 2819.3800 1035.7500 2820.0000 ;
      RECT 1028.0500 2819.3800 1031.7500 2820.0000 ;
      RECT 1024.0500 2819.3800 1027.7500 2820.0000 ;
      RECT 1020.0500 2819.3800 1023.7500 2820.0000 ;
      RECT 1016.0500 2819.3800 1019.7500 2820.0000 ;
      RECT 1012.0500 2819.3800 1015.7500 2820.0000 ;
      RECT 1008.0500 2819.3800 1011.7500 2820.0000 ;
      RECT 1004.0500 2819.3800 1007.7500 2820.0000 ;
      RECT 1000.0500 2819.3800 1003.7500 2820.0000 ;
      RECT 996.0500 2819.3800 999.7500 2820.0000 ;
      RECT 992.0500 2819.3800 995.7500 2820.0000 ;
      RECT 988.0500 2819.3800 991.7500 2820.0000 ;
      RECT 984.0500 2819.3800 987.7500 2820.0000 ;
      RECT 980.0500 2819.3800 983.7500 2820.0000 ;
      RECT 976.0500 2819.3800 979.7500 2820.0000 ;
      RECT 972.0500 2819.3800 975.7500 2820.0000 ;
      RECT 968.0500 2819.3800 971.7500 2820.0000 ;
      RECT 964.0500 2819.3800 967.7500 2820.0000 ;
      RECT 960.0500 2819.3800 963.7500 2820.0000 ;
      RECT 956.0500 2819.3800 959.7500 2820.0000 ;
      RECT 952.0500 2819.3800 955.7500 2820.0000 ;
      RECT 948.0500 2819.3800 951.7500 2820.0000 ;
      RECT 944.0500 2819.3800 947.7500 2820.0000 ;
      RECT 940.0500 2819.3800 943.7500 2820.0000 ;
      RECT 936.0500 2819.3800 939.7500 2820.0000 ;
      RECT 932.0500 2819.3800 935.7500 2820.0000 ;
      RECT 928.0500 2819.3800 931.7500 2820.0000 ;
      RECT 924.0500 2819.3800 927.7500 2820.0000 ;
      RECT 920.0500 2819.3800 923.7500 2820.0000 ;
      RECT 916.0500 2819.3800 919.7500 2820.0000 ;
      RECT 912.0500 2819.3800 915.7500 2820.0000 ;
      RECT 908.0500 2819.3800 911.7500 2820.0000 ;
      RECT 904.0500 2819.3800 907.7500 2820.0000 ;
      RECT 900.0500 2819.3800 903.7500 2820.0000 ;
      RECT 896.0500 2819.3800 899.7500 2820.0000 ;
      RECT 892.0500 2819.3800 895.7500 2820.0000 ;
      RECT 888.0500 2819.3800 891.7500 2820.0000 ;
      RECT 884.0500 2819.3800 887.7500 2820.0000 ;
      RECT 880.0500 2819.3800 883.7500 2820.0000 ;
      RECT 876.0500 2819.3800 879.7500 2820.0000 ;
      RECT 872.0500 2819.3800 875.7500 2820.0000 ;
      RECT 868.0500 2819.3800 871.7500 2820.0000 ;
      RECT 864.0500 2819.3800 867.7500 2820.0000 ;
      RECT 860.0500 2819.3800 863.7500 2820.0000 ;
      RECT 856.0500 2819.3800 859.7500 2820.0000 ;
      RECT 852.0500 2819.3800 855.7500 2820.0000 ;
      RECT 848.0500 2819.3800 851.7500 2820.0000 ;
      RECT 844.0500 2819.3800 847.7500 2820.0000 ;
      RECT 840.0500 2819.3800 843.7500 2820.0000 ;
      RECT 836.0500 2819.3800 839.7500 2820.0000 ;
      RECT 832.0500 2819.3800 835.7500 2820.0000 ;
      RECT 828.0500 2819.3800 831.7500 2820.0000 ;
      RECT 824.0500 2819.3800 827.7500 2820.0000 ;
      RECT 820.0500 2819.3800 823.7500 2820.0000 ;
      RECT 816.0500 2819.3800 819.7500 2820.0000 ;
      RECT 812.0500 2819.3800 815.7500 2820.0000 ;
      RECT 808.0500 2819.3800 811.7500 2820.0000 ;
      RECT 804.0500 2819.3800 807.7500 2820.0000 ;
      RECT 800.0500 2819.3800 803.7500 2820.0000 ;
      RECT 796.0500 2819.3800 799.7500 2820.0000 ;
      RECT 792.0500 2819.3800 795.7500 2820.0000 ;
      RECT 788.0500 2819.3800 791.7500 2820.0000 ;
      RECT 784.0500 2819.3800 787.7500 2820.0000 ;
      RECT 780.0500 2819.3800 783.7500 2820.0000 ;
      RECT 776.0500 2819.3800 779.7500 2820.0000 ;
      RECT 772.0500 2819.3800 775.7500 2820.0000 ;
      RECT 768.0500 2819.3800 771.7500 2820.0000 ;
      RECT 764.0500 2819.3800 767.7500 2820.0000 ;
      RECT 760.0500 2819.3800 763.7500 2820.0000 ;
      RECT 756.0500 2819.3800 759.7500 2820.0000 ;
      RECT 752.0500 2819.3800 755.7500 2820.0000 ;
      RECT 748.0500 2819.3800 751.7500 2820.0000 ;
      RECT 744.0500 2819.3800 747.7500 2820.0000 ;
      RECT 740.0500 2819.3800 743.7500 2820.0000 ;
      RECT 736.0500 2819.3800 739.7500 2820.0000 ;
      RECT 732.0500 2819.3800 735.7500 2820.0000 ;
      RECT 728.0500 2819.3800 731.7500 2820.0000 ;
      RECT 724.0500 2819.3800 727.7500 2820.0000 ;
      RECT 720.0500 2819.3800 723.7500 2820.0000 ;
      RECT 716.0500 2819.3800 719.7500 2820.0000 ;
      RECT 712.0500 2819.3800 715.7500 2820.0000 ;
      RECT 708.0500 2819.3800 711.7500 2820.0000 ;
      RECT 704.0500 2819.3800 707.7500 2820.0000 ;
      RECT 700.0500 2819.3800 703.7500 2820.0000 ;
      RECT 696.0500 2819.3800 699.7500 2820.0000 ;
      RECT 692.0500 2819.3800 695.7500 2820.0000 ;
      RECT 688.0500 2819.3800 691.7500 2820.0000 ;
      RECT 684.0500 2819.3800 687.7500 2820.0000 ;
      RECT 680.0500 2819.3800 683.7500 2820.0000 ;
      RECT 676.0500 2819.3800 679.7500 2820.0000 ;
      RECT 672.0500 2819.3800 675.7500 2820.0000 ;
      RECT 668.0500 2819.3800 671.7500 2820.0000 ;
      RECT 664.0500 2819.3800 667.7500 2820.0000 ;
      RECT 660.0500 2819.3800 663.7500 2820.0000 ;
      RECT 656.0500 2819.3800 659.7500 2820.0000 ;
      RECT 652.0500 2819.3800 655.7500 2820.0000 ;
      RECT 648.0500 2819.3800 651.7500 2820.0000 ;
      RECT 644.0500 2819.3800 647.7500 2820.0000 ;
      RECT 640.0500 2819.3800 643.7500 2820.0000 ;
      RECT 636.0500 2819.3800 639.7500 2820.0000 ;
      RECT 632.0500 2819.3800 635.7500 2820.0000 ;
      RECT 628.0500 2819.3800 631.7500 2820.0000 ;
      RECT 624.0500 2819.3800 627.7500 2820.0000 ;
      RECT 620.0500 2819.3800 623.7500 2820.0000 ;
      RECT 616.0500 2819.3800 619.7500 2820.0000 ;
      RECT 612.0500 2819.3800 615.7500 2820.0000 ;
      RECT 608.0500 2819.3800 611.7500 2820.0000 ;
      RECT 604.0500 2819.3800 607.7500 2820.0000 ;
      RECT 600.0500 2819.3800 603.7500 2820.0000 ;
      RECT 596.0500 2819.3800 599.7500 2820.0000 ;
      RECT 592.0500 2819.3800 595.7500 2820.0000 ;
      RECT 588.0500 2819.3800 591.7500 2820.0000 ;
      RECT 584.0500 2819.3800 587.7500 2820.0000 ;
      RECT 580.0500 2819.3800 583.7500 2820.0000 ;
      RECT 576.0500 2819.3800 579.7500 2820.0000 ;
      RECT 572.0500 2819.3800 575.7500 2820.0000 ;
      RECT 568.0500 2819.3800 571.7500 2820.0000 ;
      RECT 564.0500 2819.3800 567.7500 2820.0000 ;
      RECT 560.0500 2819.3800 563.7500 2820.0000 ;
      RECT 556.0500 2819.3800 559.7500 2820.0000 ;
      RECT 552.0500 2819.3800 555.7500 2820.0000 ;
      RECT 548.0500 2819.3800 551.7500 2820.0000 ;
      RECT 544.0500 2819.3800 547.7500 2820.0000 ;
      RECT 540.0500 2819.3800 543.7500 2820.0000 ;
      RECT 536.0500 2819.3800 539.7500 2820.0000 ;
      RECT 532.0500 2819.3800 535.7500 2820.0000 ;
      RECT 528.0500 2819.3800 531.7500 2820.0000 ;
      RECT 524.0500 2819.3800 527.7500 2820.0000 ;
      RECT 520.0500 2819.3800 523.7500 2820.0000 ;
      RECT 516.0500 2819.3800 519.7500 2820.0000 ;
      RECT 512.0500 2819.3800 515.7500 2820.0000 ;
      RECT 508.0500 2819.3800 511.7500 2820.0000 ;
      RECT 504.0500 2819.3800 507.7500 2820.0000 ;
      RECT 500.0500 2819.3800 503.7500 2820.0000 ;
      RECT 496.0500 2819.3800 499.7500 2820.0000 ;
      RECT 492.0500 2819.3800 495.7500 2820.0000 ;
      RECT 488.0500 2819.3800 491.7500 2820.0000 ;
      RECT 484.0500 2819.3800 487.7500 2820.0000 ;
      RECT 480.0500 2819.3800 483.7500 2820.0000 ;
      RECT 476.0500 2819.3800 479.7500 2820.0000 ;
      RECT 472.0500 2819.3800 475.7500 2820.0000 ;
      RECT 468.0500 2819.3800 471.7500 2820.0000 ;
      RECT 464.0500 2819.3800 467.7500 2820.0000 ;
      RECT 460.0500 2819.3800 463.7500 2820.0000 ;
      RECT 456.0500 2819.3800 459.7500 2820.0000 ;
      RECT 452.0500 2819.3800 455.7500 2820.0000 ;
      RECT 448.0500 2819.3800 451.7500 2820.0000 ;
      RECT 444.0500 2819.3800 447.7500 2820.0000 ;
      RECT 440.0500 2819.3800 443.7500 2820.0000 ;
      RECT 436.0500 2819.3800 439.7500 2820.0000 ;
      RECT 432.0500 2819.3800 435.7500 2820.0000 ;
      RECT 428.0500 2819.3800 431.7500 2820.0000 ;
      RECT 424.0500 2819.3800 427.7500 2820.0000 ;
      RECT 420.0500 2819.3800 423.7500 2820.0000 ;
      RECT 416.0500 2819.3800 419.7500 2820.0000 ;
      RECT 412.0500 2819.3800 415.7500 2820.0000 ;
      RECT 408.0500 2819.3800 411.7500 2820.0000 ;
      RECT 404.0500 2819.3800 407.7500 2820.0000 ;
      RECT 400.0500 2819.3800 403.7500 2820.0000 ;
      RECT 396.0500 2819.3800 399.7500 2820.0000 ;
      RECT 392.0500 2819.3800 395.7500 2820.0000 ;
      RECT 388.0500 2819.3800 391.7500 2820.0000 ;
      RECT 384.0500 2819.3800 387.7500 2820.0000 ;
      RECT 380.0500 2819.3800 383.7500 2820.0000 ;
      RECT 376.0500 2819.3800 379.7500 2820.0000 ;
      RECT 372.0500 2819.3800 375.7500 2820.0000 ;
      RECT 368.0500 2819.3800 371.7500 2820.0000 ;
      RECT 364.0500 2819.3800 367.7500 2820.0000 ;
      RECT 360.0500 2819.3800 363.7500 2820.0000 ;
      RECT 356.0500 2819.3800 359.7500 2820.0000 ;
      RECT 352.0500 2819.3800 355.7500 2820.0000 ;
      RECT 348.0500 2819.3800 351.7500 2820.0000 ;
      RECT 344.0500 2819.3800 347.7500 2820.0000 ;
      RECT 340.0500 2819.3800 343.7500 2820.0000 ;
      RECT 336.0500 2819.3800 339.7500 2820.0000 ;
      RECT 332.0500 2819.3800 335.7500 2820.0000 ;
      RECT 328.0500 2819.3800 331.7500 2820.0000 ;
      RECT 324.0500 2819.3800 327.7500 2820.0000 ;
      RECT 320.0500 2819.3800 323.7500 2820.0000 ;
      RECT 316.0500 2819.3800 319.7500 2820.0000 ;
      RECT 312.0500 2819.3800 315.7500 2820.0000 ;
      RECT 308.0500 2819.3800 311.7500 2820.0000 ;
      RECT 304.0500 2819.3800 307.7500 2820.0000 ;
      RECT 300.0500 2819.3800 303.7500 2820.0000 ;
      RECT 296.0500 2819.3800 299.7500 2820.0000 ;
      RECT 292.0500 2819.3800 295.7500 2820.0000 ;
      RECT 288.0500 2819.3800 291.7500 2820.0000 ;
      RECT 284.0500 2819.3800 287.7500 2820.0000 ;
      RECT 280.0500 2819.3800 283.7500 2820.0000 ;
      RECT 276.0500 2819.3800 279.7500 2820.0000 ;
      RECT 272.0500 2819.3800 275.7500 2820.0000 ;
      RECT 268.0500 2819.3800 271.7500 2820.0000 ;
      RECT 264.0500 2819.3800 267.7500 2820.0000 ;
      RECT 260.0500 2819.3800 263.7500 2820.0000 ;
      RECT 256.0500 2819.3800 259.7500 2820.0000 ;
      RECT 252.0500 2819.3800 255.7500 2820.0000 ;
      RECT 248.0500 2819.3800 251.7500 2820.0000 ;
      RECT 244.0500 2819.3800 247.7500 2820.0000 ;
      RECT 240.0500 2819.3800 243.7500 2820.0000 ;
      RECT 236.0500 2819.3800 239.7500 2820.0000 ;
      RECT 232.0500 2819.3800 235.7500 2820.0000 ;
      RECT 228.0500 2819.3800 231.7500 2820.0000 ;
      RECT 224.0500 2819.3800 227.7500 2820.0000 ;
      RECT 220.0500 2819.3800 223.7500 2820.0000 ;
      RECT 216.0500 2819.3800 219.7500 2820.0000 ;
      RECT 212.0500 2819.3800 215.7500 2820.0000 ;
      RECT 208.0500 2819.3800 211.7500 2820.0000 ;
      RECT 204.0500 2819.3800 207.7500 2820.0000 ;
      RECT 200.0500 2819.3800 203.7500 2820.0000 ;
      RECT 196.0500 2819.3800 199.7500 2820.0000 ;
      RECT 192.0500 2819.3800 195.7500 2820.0000 ;
      RECT 188.0500 2819.3800 191.7500 2820.0000 ;
      RECT 184.0500 2819.3800 187.7500 2820.0000 ;
      RECT 180.0500 2819.3800 183.7500 2820.0000 ;
      RECT 176.0500 2819.3800 179.7500 2820.0000 ;
      RECT 172.0500 2819.3800 175.7500 2820.0000 ;
      RECT 168.0500 2819.3800 171.7500 2820.0000 ;
      RECT 164.0500 2819.3800 167.7500 2820.0000 ;
      RECT 160.0500 2819.3800 163.7500 2820.0000 ;
      RECT 156.0500 2819.3800 159.7500 2820.0000 ;
      RECT 152.0500 2819.3800 155.7500 2820.0000 ;
      RECT 148.0500 2819.3800 151.7500 2820.0000 ;
      RECT 144.0500 2819.3800 147.7500 2820.0000 ;
      RECT 140.0500 2819.3800 143.7500 2820.0000 ;
      RECT 136.0500 2819.3800 139.7500 2820.0000 ;
      RECT 132.0500 2819.3800 135.7500 2820.0000 ;
      RECT 128.0500 2819.3800 131.7500 2820.0000 ;
      RECT 124.0500 2819.3800 127.7500 2820.0000 ;
      RECT 120.0500 2819.3800 123.7500 2820.0000 ;
      RECT 116.0500 2819.3800 119.7500 2820.0000 ;
      RECT 112.0500 2819.3800 115.7500 2820.0000 ;
      RECT 108.0500 2819.3800 111.7500 2820.0000 ;
      RECT 104.0500 2819.3800 107.7500 2820.0000 ;
      RECT 100.0500 2819.3800 103.7500 2820.0000 ;
      RECT 96.0500 2819.3800 99.7500 2820.0000 ;
      RECT 92.0500 2819.3800 95.7500 2820.0000 ;
      RECT 88.0500 2819.3800 91.7500 2820.0000 ;
      RECT 84.0500 2819.3800 87.7500 2820.0000 ;
      RECT 80.0500 2819.3800 83.7500 2820.0000 ;
      RECT 76.0500 2819.3800 79.7500 2820.0000 ;
      RECT 72.0500 2819.3800 75.7500 2820.0000 ;
      RECT 0.0000 2819.3800 71.7500 2820.0000 ;
      RECT 0.0000 0.6200 1420.0000 2819.3800 ;
      RECT 1006.2500 0.0000 1420.0000 0.6200 ;
      RECT 1002.2500 0.0000 1005.9500 0.6200 ;
      RECT 998.2500 0.0000 1001.9500 0.6200 ;
      RECT 994.2500 0.0000 997.9500 0.6200 ;
      RECT 990.2500 0.0000 993.9500 0.6200 ;
      RECT 986.2500 0.0000 989.9500 0.6200 ;
      RECT 982.2500 0.0000 985.9500 0.6200 ;
      RECT 978.2500 0.0000 981.9500 0.6200 ;
      RECT 974.2500 0.0000 977.9500 0.6200 ;
      RECT 970.2500 0.0000 973.9500 0.6200 ;
      RECT 966.2500 0.0000 969.9500 0.6200 ;
      RECT 962.2500 0.0000 965.9500 0.6200 ;
      RECT 958.2500 0.0000 961.9500 0.6200 ;
      RECT 954.2500 0.0000 957.9500 0.6200 ;
      RECT 950.2500 0.0000 953.9500 0.6200 ;
      RECT 946.2500 0.0000 949.9500 0.6200 ;
      RECT 942.2500 0.0000 945.9500 0.6200 ;
      RECT 938.2500 0.0000 941.9500 0.6200 ;
      RECT 934.2500 0.0000 937.9500 0.6200 ;
      RECT 930.2500 0.0000 933.9500 0.6200 ;
      RECT 926.2500 0.0000 929.9500 0.6200 ;
      RECT 922.2500 0.0000 925.9500 0.6200 ;
      RECT 918.2500 0.0000 921.9500 0.6200 ;
      RECT 914.2500 0.0000 917.9500 0.6200 ;
      RECT 910.2500 0.0000 913.9500 0.6200 ;
      RECT 906.2500 0.0000 909.9500 0.6200 ;
      RECT 902.2500 0.0000 905.9500 0.6200 ;
      RECT 898.2500 0.0000 901.9500 0.6200 ;
      RECT 894.2500 0.0000 897.9500 0.6200 ;
      RECT 890.2500 0.0000 893.9500 0.6200 ;
      RECT 886.2500 0.0000 889.9500 0.6200 ;
      RECT 882.2500 0.0000 885.9500 0.6200 ;
      RECT 878.2500 0.0000 881.9500 0.6200 ;
      RECT 874.2500 0.0000 877.9500 0.6200 ;
      RECT 870.2500 0.0000 873.9500 0.6200 ;
      RECT 866.2500 0.0000 869.9500 0.6200 ;
      RECT 862.2500 0.0000 865.9500 0.6200 ;
      RECT 858.2500 0.0000 861.9500 0.6200 ;
      RECT 854.2500 0.0000 857.9500 0.6200 ;
      RECT 850.2500 0.0000 853.9500 0.6200 ;
      RECT 846.2500 0.0000 849.9500 0.6200 ;
      RECT 842.2500 0.0000 845.9500 0.6200 ;
      RECT 838.2500 0.0000 841.9500 0.6200 ;
      RECT 834.2500 0.0000 837.9500 0.6200 ;
      RECT 830.2500 0.0000 833.9500 0.6200 ;
      RECT 826.2500 0.0000 829.9500 0.6200 ;
      RECT 822.2500 0.0000 825.9500 0.6200 ;
      RECT 818.2500 0.0000 821.9500 0.6200 ;
      RECT 814.2500 0.0000 817.9500 0.6200 ;
      RECT 810.2500 0.0000 813.9500 0.6200 ;
      RECT 806.2500 0.0000 809.9500 0.6200 ;
      RECT 802.2500 0.0000 805.9500 0.6200 ;
      RECT 798.2500 0.0000 801.9500 0.6200 ;
      RECT 794.2500 0.0000 797.9500 0.6200 ;
      RECT 790.2500 0.0000 793.9500 0.6200 ;
      RECT 786.2500 0.0000 789.9500 0.6200 ;
      RECT 782.2500 0.0000 785.9500 0.6200 ;
      RECT 778.2500 0.0000 781.9500 0.6200 ;
      RECT 774.2500 0.0000 777.9500 0.6200 ;
      RECT 770.2500 0.0000 773.9500 0.6200 ;
      RECT 766.2500 0.0000 769.9500 0.6200 ;
      RECT 762.2500 0.0000 765.9500 0.6200 ;
      RECT 758.2500 0.0000 761.9500 0.6200 ;
      RECT 754.2500 0.0000 757.9500 0.6200 ;
      RECT 750.2500 0.0000 753.9500 0.6200 ;
      RECT 746.2500 0.0000 749.9500 0.6200 ;
      RECT 742.2500 0.0000 745.9500 0.6200 ;
      RECT 738.2500 0.0000 741.9500 0.6200 ;
      RECT 734.2500 0.0000 737.9500 0.6200 ;
      RECT 730.2500 0.0000 733.9500 0.6200 ;
      RECT 726.2500 0.0000 729.9500 0.6200 ;
      RECT 722.2500 0.0000 725.9500 0.6200 ;
      RECT 718.2500 0.0000 721.9500 0.6200 ;
      RECT 714.2500 0.0000 717.9500 0.6200 ;
      RECT 710.2500 0.0000 713.9500 0.6200 ;
      RECT 706.2500 0.0000 709.9500 0.6200 ;
      RECT 702.2500 0.0000 705.9500 0.6200 ;
      RECT 698.2500 0.0000 701.9500 0.6200 ;
      RECT 694.2500 0.0000 697.9500 0.6200 ;
      RECT 690.2500 0.0000 693.9500 0.6200 ;
      RECT 686.2500 0.0000 689.9500 0.6200 ;
      RECT 682.2500 0.0000 685.9500 0.6200 ;
      RECT 678.2500 0.0000 681.9500 0.6200 ;
      RECT 674.2500 0.0000 677.9500 0.6200 ;
      RECT 670.2500 0.0000 673.9500 0.6200 ;
      RECT 666.2500 0.0000 669.9500 0.6200 ;
      RECT 662.2500 0.0000 665.9500 0.6200 ;
      RECT 658.2500 0.0000 661.9500 0.6200 ;
      RECT 654.2500 0.0000 657.9500 0.6200 ;
      RECT 650.2500 0.0000 653.9500 0.6200 ;
      RECT 646.2500 0.0000 649.9500 0.6200 ;
      RECT 642.2500 0.0000 645.9500 0.6200 ;
      RECT 638.2500 0.0000 641.9500 0.6200 ;
      RECT 634.2500 0.0000 637.9500 0.6200 ;
      RECT 630.2500 0.0000 633.9500 0.6200 ;
      RECT 626.2500 0.0000 629.9500 0.6200 ;
      RECT 622.2500 0.0000 625.9500 0.6200 ;
      RECT 618.2500 0.0000 621.9500 0.6200 ;
      RECT 614.2500 0.0000 617.9500 0.6200 ;
      RECT 610.2500 0.0000 613.9500 0.6200 ;
      RECT 606.2500 0.0000 609.9500 0.6200 ;
      RECT 602.2500 0.0000 605.9500 0.6200 ;
      RECT 598.2500 0.0000 601.9500 0.6200 ;
      RECT 594.2500 0.0000 597.9500 0.6200 ;
      RECT 590.2500 0.0000 593.9500 0.6200 ;
      RECT 586.2500 0.0000 589.9500 0.6200 ;
      RECT 582.2500 0.0000 585.9500 0.6200 ;
      RECT 578.2500 0.0000 581.9500 0.6200 ;
      RECT 574.2500 0.0000 577.9500 0.6200 ;
      RECT 570.2500 0.0000 573.9500 0.6200 ;
      RECT 566.2500 0.0000 569.9500 0.6200 ;
      RECT 562.2500 0.0000 565.9500 0.6200 ;
      RECT 558.2500 0.0000 561.9500 0.6200 ;
      RECT 554.2500 0.0000 557.9500 0.6200 ;
      RECT 550.2500 0.0000 553.9500 0.6200 ;
      RECT 546.2500 0.0000 549.9500 0.6200 ;
      RECT 542.2500 0.0000 545.9500 0.6200 ;
      RECT 538.2500 0.0000 541.9500 0.6200 ;
      RECT 534.2500 0.0000 537.9500 0.6200 ;
      RECT 530.2500 0.0000 533.9500 0.6200 ;
      RECT 526.2500 0.0000 529.9500 0.6200 ;
      RECT 522.2500 0.0000 525.9500 0.6200 ;
      RECT 518.2500 0.0000 521.9500 0.6200 ;
      RECT 514.2500 0.0000 517.9500 0.6200 ;
      RECT 510.2500 0.0000 513.9500 0.6200 ;
      RECT 506.2500 0.0000 509.9500 0.6200 ;
      RECT 502.2500 0.0000 505.9500 0.6200 ;
      RECT 498.2500 0.0000 501.9500 0.6200 ;
      RECT 494.2500 0.0000 497.9500 0.6200 ;
      RECT 490.2500 0.0000 493.9500 0.6200 ;
      RECT 486.2500 0.0000 489.9500 0.6200 ;
      RECT 482.2500 0.0000 485.9500 0.6200 ;
      RECT 478.2500 0.0000 481.9500 0.6200 ;
      RECT 474.2500 0.0000 477.9500 0.6200 ;
      RECT 470.2500 0.0000 473.9500 0.6200 ;
      RECT 466.2500 0.0000 469.9500 0.6200 ;
      RECT 462.2500 0.0000 465.9500 0.6200 ;
      RECT 458.2500 0.0000 461.9500 0.6200 ;
      RECT 454.2500 0.0000 457.9500 0.6200 ;
      RECT 450.2500 0.0000 453.9500 0.6200 ;
      RECT 446.2500 0.0000 449.9500 0.6200 ;
      RECT 442.2500 0.0000 445.9500 0.6200 ;
      RECT 438.2500 0.0000 441.9500 0.6200 ;
      RECT 434.2500 0.0000 437.9500 0.6200 ;
      RECT 430.2500 0.0000 433.9500 0.6200 ;
      RECT 426.2500 0.0000 429.9500 0.6200 ;
      RECT 422.2500 0.0000 425.9500 0.6200 ;
      RECT 418.2500 0.0000 421.9500 0.6200 ;
      RECT 414.2500 0.0000 417.9500 0.6200 ;
      RECT 0.0000 0.0000 413.9500 0.6200 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 1420.0000 2820.0000 ;
  END
END fullchip

END LIBRARY
