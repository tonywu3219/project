/home/linux/ieng6/ee260bwi25/zuy001/project/project/project_p3/pnr_core/subckt/sram_w16_64b.lef