##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sun Mar 16 13:55:00 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 540.0000 BY 540.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 267.2550 539.5300 267.3450 540.0000 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 389.7500 0.5200 389.8500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 386.7500 0.5200 386.8500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 383.7500 0.5200 383.8500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 380.7500 0.5200 380.8500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 377.7500 0.5200 377.8500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 374.7500 0.5200 374.8500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 371.7500 0.5200 371.8500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 368.7500 0.5200 368.8500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 365.7500 0.5200 365.8500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 362.7500 0.5200 362.8500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 359.7500 0.5200 359.8500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 356.7500 0.5200 356.8500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 353.7500 0.5200 353.8500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 350.7500 0.5200 350.8500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 347.7500 0.5200 347.8500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 344.7500 0.5200 344.8500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 341.7500 0.5200 341.8500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 338.7500 0.5200 338.8500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 335.7500 0.5200 335.8500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 332.7500 0.5200 332.8500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 329.7500 0.5200 329.8500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 326.7500 0.5200 326.8500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 323.7500 0.5200 323.8500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 320.7500 0.5200 320.8500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 317.7500 0.5200 317.8500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 314.7500 0.5200 314.8500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 311.7500 0.5200 311.8500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 308.7500 0.5200 308.8500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 305.7500 0.5200 305.8500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 302.7500 0.5200 302.8500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 299.7500 0.5200 299.8500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 296.7500 0.5200 296.8500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 293.7500 0.5200 293.8500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 290.7500 0.5200 290.8500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 287.7500 0.5200 287.8500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 284.7500 0.5200 284.8500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 281.7500 0.5200 281.8500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 278.7500 0.5200 278.8500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 275.7500 0.5200 275.8500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 272.7500 0.5200 272.8500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 269.7500 0.5200 269.8500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 266.7500 0.5200 266.8500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 263.7500 0.5200 263.8500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 260.7500 0.5200 260.8500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 257.7500 0.5200 257.8500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 254.7500 0.5200 254.8500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 251.7500 0.5200 251.8500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 248.7500 0.5200 248.8500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 245.7500 0.5200 245.8500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 242.7500 0.5200 242.8500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 239.7500 0.5200 239.8500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 236.7500 0.5200 236.8500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 233.7500 0.5200 233.8500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 230.7500 0.5200 230.8500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 227.7500 0.5200 227.8500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 224.7500 0.5200 224.8500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 221.7500 0.5200 221.8500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 218.7500 0.5200 218.8500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 215.7500 0.5200 215.8500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 212.7500 0.5200 212.8500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 209.7500 0.5200 209.8500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 206.7500 0.5200 206.8500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 203.7500 0.5200 203.8500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 200.7500 0.5200 200.8500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 428.8550 0.0000 428.9450 0.4700 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 426.8550 0.0000 426.9450 0.4700 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 424.8550 0.0000 424.9450 0.4700 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 422.8550 0.0000 422.9450 0.4700 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 420.8550 0.0000 420.9450 0.4700 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 418.8550 0.0000 418.9450 0.4700 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 416.8550 0.0000 416.9450 0.4700 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 414.8550 0.0000 414.9450 0.4700 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 412.8550 0.0000 412.9450 0.4700 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 410.8550 0.0000 410.9450 0.4700 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 408.8550 0.0000 408.9450 0.4700 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 406.8550 0.0000 406.9450 0.4700 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 404.8550 0.0000 404.9450 0.4700 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 402.8550 0.0000 402.9450 0.4700 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 400.8550 0.0000 400.9450 0.4700 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 398.8550 0.0000 398.9450 0.4700 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 396.8550 0.0000 396.9450 0.4700 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 394.8550 0.0000 394.9450 0.4700 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 392.8550 0.0000 392.9450 0.4700 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 390.8550 0.0000 390.9450 0.4700 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 388.8550 0.0000 388.9450 0.4700 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 386.8550 0.0000 386.9450 0.4700 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 384.8550 0.0000 384.9450 0.4700 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 382.8550 0.0000 382.9450 0.4700 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 380.8550 0.0000 380.9450 0.4700 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 378.8550 0.0000 378.9450 0.4700 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 376.8550 0.0000 376.9450 0.4700 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 374.8550 0.0000 374.9450 0.4700 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 372.8550 0.0000 372.9450 0.4700 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 370.8550 0.0000 370.9450 0.4700 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 368.8550 0.0000 368.9450 0.4700 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 366.8550 0.0000 366.9450 0.4700 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 364.8550 0.0000 364.9450 0.4700 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 362.8550 0.0000 362.9450 0.4700 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 360.8550 0.0000 360.9450 0.4700 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 358.8550 0.0000 358.9450 0.4700 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 356.8550 0.0000 356.9450 0.4700 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 354.8550 0.0000 354.9450 0.4700 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 352.8550 0.0000 352.9450 0.4700 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 350.8550 0.0000 350.9450 0.4700 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 348.8550 0.0000 348.9450 0.4700 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 346.8550 0.0000 346.9450 0.4700 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 344.8550 0.0000 344.9450 0.4700 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 342.8550 0.0000 342.9450 0.4700 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 340.8550 0.0000 340.9450 0.4700 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 338.8550 0.0000 338.9450 0.4700 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 336.8550 0.0000 336.9450 0.4700 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 334.8550 0.0000 334.9450 0.4700 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 332.8550 0.0000 332.9450 0.4700 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 330.8550 0.0000 330.9450 0.4700 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 328.8550 0.0000 328.9450 0.4700 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 326.8550 0.0000 326.9450 0.4700 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 324.8550 0.0000 324.9450 0.4700 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 322.8550 0.0000 322.9450 0.4700 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 320.8550 0.0000 320.9450 0.4700 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 318.8550 0.0000 318.9450 0.4700 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 316.8550 0.0000 316.9450 0.4700 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 314.8550 0.0000 314.9450 0.4700 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 312.8550 0.0000 312.9450 0.4700 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 310.8550 0.0000 310.9450 0.4700 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 308.8550 0.0000 308.9450 0.4700 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 306.8550 0.0000 306.9450 0.4700 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 304.8550 0.0000 304.9450 0.4700 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 302.8550 0.0000 302.9450 0.4700 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 300.8550 0.0000 300.9450 0.4700 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 298.8550 0.0000 298.9450 0.4700 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 296.8550 0.0000 296.9450 0.4700 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 294.8550 0.0000 294.9450 0.4700 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 292.8550 0.0000 292.9450 0.4700 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 290.8550 0.0000 290.9450 0.4700 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 288.8550 0.0000 288.9450 0.4700 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 286.8550 0.0000 286.9450 0.4700 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 284.8550 0.0000 284.9450 0.4700 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 282.8550 0.0000 282.9450 0.4700 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 280.8550 0.0000 280.9450 0.4700 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 278.8550 0.0000 278.9450 0.4700 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 276.8550 0.0000 276.9450 0.4700 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 274.8550 0.0000 274.9450 0.4700 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 272.8550 0.0000 272.9450 0.4700 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 270.8550 0.0000 270.9450 0.4700 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 268.8550 0.0000 268.9450 0.4700 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 266.8550 0.0000 266.9450 0.4700 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 264.8550 0.0000 264.9450 0.4700 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 262.8550 0.0000 262.9450 0.4700 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 260.8550 0.0000 260.9450 0.4700 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 258.8550 0.0000 258.9450 0.4700 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 256.8550 0.0000 256.9450 0.4700 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 254.8550 0.0000 254.9450 0.4700 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 252.8550 0.0000 252.9450 0.4700 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 250.8550 0.0000 250.9450 0.4700 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 248.8550 0.0000 248.9450 0.4700 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 246.8550 0.0000 246.9450 0.4700 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 244.8550 0.0000 244.9450 0.4700 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 242.8550 0.0000 242.9450 0.4700 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 240.8550 0.0000 240.9450 0.4700 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 238.8550 0.0000 238.9450 0.4700 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 236.8550 0.0000 236.9450 0.4700 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 234.8550 0.0000 234.9450 0.4700 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 232.8550 0.0000 232.9450 0.4700 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 230.8550 0.0000 230.9450 0.4700 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 228.8550 0.0000 228.9450 0.4700 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 226.8550 0.0000 226.9450 0.4700 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 224.8550 0.0000 224.9450 0.4700 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 222.8550 0.0000 222.9450 0.4700 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 220.8550 0.0000 220.9450 0.4700 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 218.8550 0.0000 218.9450 0.4700 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 216.8550 0.0000 216.9450 0.4700 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 214.8550 0.0000 214.9450 0.4700 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 212.8550 0.0000 212.9450 0.4700 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 210.8550 0.0000 210.9450 0.4700 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 208.8550 0.0000 208.9450 0.4700 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 206.8550 0.0000 206.9450 0.4700 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 204.8550 0.0000 204.9450 0.4700 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 202.8550 0.0000 202.9450 0.4700 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 200.8550 0.0000 200.9450 0.4700 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 198.8550 0.0000 198.9450 0.4700 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 196.8550 0.0000 196.9450 0.4700 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 194.8550 0.0000 194.9450 0.4700 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 192.8550 0.0000 192.9450 0.4700 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 190.8550 0.0000 190.9450 0.4700 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 188.8550 0.0000 188.9450 0.4700 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 186.8550 0.0000 186.9450 0.4700 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 184.8550 0.0000 184.9450 0.4700 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 182.8550 0.0000 182.9450 0.4700 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 180.8550 0.0000 180.9450 0.4700 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 178.8550 0.0000 178.9450 0.4700 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 176.8550 0.0000 176.9450 0.4700 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 174.8550 0.0000 174.9450 0.4700 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 172.8550 0.0000 172.9450 0.4700 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 170.8550 0.0000 170.9450 0.4700 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 168.8550 0.0000 168.9450 0.4700 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 166.8550 0.0000 166.9450 0.4700 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 164.8550 0.0000 164.9450 0.4700 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 162.8550 0.0000 162.9450 0.4700 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 160.8550 0.0000 160.9450 0.4700 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 158.8550 0.0000 158.9450 0.4700 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 156.8550 0.0000 156.9450 0.4700 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 154.8550 0.0000 154.9450 0.4700 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 152.8550 0.0000 152.9450 0.4700 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 150.8550 0.0000 150.9450 0.4700 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 148.8550 0.0000 148.9450 0.4700 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 146.8550 0.0000 146.9450 0.4700 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 144.8550 0.0000 144.9450 0.4700 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 142.8550 0.0000 142.9450 0.4700 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 140.8550 0.0000 140.9450 0.4700 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 138.8550 0.0000 138.9450 0.4700 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 136.8550 0.0000 136.9450 0.4700 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 134.8550 0.0000 134.9450 0.4700 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 132.8550 0.0000 132.9450 0.4700 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 130.8550 0.0000 130.9450 0.4700 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 128.8550 0.0000 128.9450 0.4700 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 126.8550 0.0000 126.9450 0.4700 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 124.8550 0.0000 124.9450 0.4700 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 122.8550 0.0000 122.9450 0.4700 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 120.8550 0.0000 120.9450 0.4700 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 118.8550 0.0000 118.9450 0.4700 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 116.8550 0.0000 116.9450 0.4700 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 114.8550 0.0000 114.9450 0.4700 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 112.8550 0.0000 112.9450 0.4700 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 110.8550 0.0000 110.9450 0.4700 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 197.7500 0.5200 197.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 194.7500 0.5200 194.8500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 191.7500 0.5200 191.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 188.7500 0.5200 188.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 185.7500 0.5200 185.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 182.7500 0.5200 182.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 179.7500 0.5200 179.8500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 176.7500 0.5200 176.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 173.7500 0.5200 173.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 170.7500 0.5200 170.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 167.7500 0.5200 167.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 164.7500 0.5200 164.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 161.7500 0.5200 161.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 158.7500 0.5200 158.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 155.7500 0.5200 155.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 152.7500 0.5200 152.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 149.7500 0.5200 149.8500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 272.2550 539.5300 272.3450 540.0000 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 272.5050 539.3700 540.0000 540.0000 ;
      RECT 267.5050 539.3700 272.0950 540.0000 ;
      RECT 0.0000 539.3700 267.0950 540.0000 ;
      RECT 0.0000 0.6300 540.0000 539.3700 ;
      RECT 429.1050 0.0000 540.0000 0.6300 ;
      RECT 427.1050 0.0000 428.6950 0.6300 ;
      RECT 425.1050 0.0000 426.6950 0.6300 ;
      RECT 423.1050 0.0000 424.6950 0.6300 ;
      RECT 421.1050 0.0000 422.6950 0.6300 ;
      RECT 419.1050 0.0000 420.6950 0.6300 ;
      RECT 417.1050 0.0000 418.6950 0.6300 ;
      RECT 415.1050 0.0000 416.6950 0.6300 ;
      RECT 413.1050 0.0000 414.6950 0.6300 ;
      RECT 411.1050 0.0000 412.6950 0.6300 ;
      RECT 409.1050 0.0000 410.6950 0.6300 ;
      RECT 407.1050 0.0000 408.6950 0.6300 ;
      RECT 405.1050 0.0000 406.6950 0.6300 ;
      RECT 403.1050 0.0000 404.6950 0.6300 ;
      RECT 401.1050 0.0000 402.6950 0.6300 ;
      RECT 399.1050 0.0000 400.6950 0.6300 ;
      RECT 397.1050 0.0000 398.6950 0.6300 ;
      RECT 395.1050 0.0000 396.6950 0.6300 ;
      RECT 393.1050 0.0000 394.6950 0.6300 ;
      RECT 391.1050 0.0000 392.6950 0.6300 ;
      RECT 389.1050 0.0000 390.6950 0.6300 ;
      RECT 387.1050 0.0000 388.6950 0.6300 ;
      RECT 385.1050 0.0000 386.6950 0.6300 ;
      RECT 383.1050 0.0000 384.6950 0.6300 ;
      RECT 381.1050 0.0000 382.6950 0.6300 ;
      RECT 379.1050 0.0000 380.6950 0.6300 ;
      RECT 377.1050 0.0000 378.6950 0.6300 ;
      RECT 375.1050 0.0000 376.6950 0.6300 ;
      RECT 373.1050 0.0000 374.6950 0.6300 ;
      RECT 371.1050 0.0000 372.6950 0.6300 ;
      RECT 369.1050 0.0000 370.6950 0.6300 ;
      RECT 367.1050 0.0000 368.6950 0.6300 ;
      RECT 365.1050 0.0000 366.6950 0.6300 ;
      RECT 363.1050 0.0000 364.6950 0.6300 ;
      RECT 361.1050 0.0000 362.6950 0.6300 ;
      RECT 359.1050 0.0000 360.6950 0.6300 ;
      RECT 357.1050 0.0000 358.6950 0.6300 ;
      RECT 355.1050 0.0000 356.6950 0.6300 ;
      RECT 353.1050 0.0000 354.6950 0.6300 ;
      RECT 351.1050 0.0000 352.6950 0.6300 ;
      RECT 349.1050 0.0000 350.6950 0.6300 ;
      RECT 347.1050 0.0000 348.6950 0.6300 ;
      RECT 345.1050 0.0000 346.6950 0.6300 ;
      RECT 343.1050 0.0000 344.6950 0.6300 ;
      RECT 341.1050 0.0000 342.6950 0.6300 ;
      RECT 339.1050 0.0000 340.6950 0.6300 ;
      RECT 337.1050 0.0000 338.6950 0.6300 ;
      RECT 335.1050 0.0000 336.6950 0.6300 ;
      RECT 333.1050 0.0000 334.6950 0.6300 ;
      RECT 331.1050 0.0000 332.6950 0.6300 ;
      RECT 329.1050 0.0000 330.6950 0.6300 ;
      RECT 327.1050 0.0000 328.6950 0.6300 ;
      RECT 325.1050 0.0000 326.6950 0.6300 ;
      RECT 323.1050 0.0000 324.6950 0.6300 ;
      RECT 321.1050 0.0000 322.6950 0.6300 ;
      RECT 319.1050 0.0000 320.6950 0.6300 ;
      RECT 317.1050 0.0000 318.6950 0.6300 ;
      RECT 315.1050 0.0000 316.6950 0.6300 ;
      RECT 313.1050 0.0000 314.6950 0.6300 ;
      RECT 311.1050 0.0000 312.6950 0.6300 ;
      RECT 309.1050 0.0000 310.6950 0.6300 ;
      RECT 307.1050 0.0000 308.6950 0.6300 ;
      RECT 305.1050 0.0000 306.6950 0.6300 ;
      RECT 303.1050 0.0000 304.6950 0.6300 ;
      RECT 301.1050 0.0000 302.6950 0.6300 ;
      RECT 299.1050 0.0000 300.6950 0.6300 ;
      RECT 297.1050 0.0000 298.6950 0.6300 ;
      RECT 295.1050 0.0000 296.6950 0.6300 ;
      RECT 293.1050 0.0000 294.6950 0.6300 ;
      RECT 291.1050 0.0000 292.6950 0.6300 ;
      RECT 289.1050 0.0000 290.6950 0.6300 ;
      RECT 287.1050 0.0000 288.6950 0.6300 ;
      RECT 285.1050 0.0000 286.6950 0.6300 ;
      RECT 283.1050 0.0000 284.6950 0.6300 ;
      RECT 281.1050 0.0000 282.6950 0.6300 ;
      RECT 279.1050 0.0000 280.6950 0.6300 ;
      RECT 277.1050 0.0000 278.6950 0.6300 ;
      RECT 275.1050 0.0000 276.6950 0.6300 ;
      RECT 273.1050 0.0000 274.6950 0.6300 ;
      RECT 271.1050 0.0000 272.6950 0.6300 ;
      RECT 269.1050 0.0000 270.6950 0.6300 ;
      RECT 267.1050 0.0000 268.6950 0.6300 ;
      RECT 265.1050 0.0000 266.6950 0.6300 ;
      RECT 263.1050 0.0000 264.6950 0.6300 ;
      RECT 261.1050 0.0000 262.6950 0.6300 ;
      RECT 259.1050 0.0000 260.6950 0.6300 ;
      RECT 257.1050 0.0000 258.6950 0.6300 ;
      RECT 255.1050 0.0000 256.6950 0.6300 ;
      RECT 253.1050 0.0000 254.6950 0.6300 ;
      RECT 251.1050 0.0000 252.6950 0.6300 ;
      RECT 249.1050 0.0000 250.6950 0.6300 ;
      RECT 247.1050 0.0000 248.6950 0.6300 ;
      RECT 245.1050 0.0000 246.6950 0.6300 ;
      RECT 243.1050 0.0000 244.6950 0.6300 ;
      RECT 241.1050 0.0000 242.6950 0.6300 ;
      RECT 239.1050 0.0000 240.6950 0.6300 ;
      RECT 237.1050 0.0000 238.6950 0.6300 ;
      RECT 235.1050 0.0000 236.6950 0.6300 ;
      RECT 233.1050 0.0000 234.6950 0.6300 ;
      RECT 231.1050 0.0000 232.6950 0.6300 ;
      RECT 229.1050 0.0000 230.6950 0.6300 ;
      RECT 227.1050 0.0000 228.6950 0.6300 ;
      RECT 225.1050 0.0000 226.6950 0.6300 ;
      RECT 223.1050 0.0000 224.6950 0.6300 ;
      RECT 221.1050 0.0000 222.6950 0.6300 ;
      RECT 219.1050 0.0000 220.6950 0.6300 ;
      RECT 217.1050 0.0000 218.6950 0.6300 ;
      RECT 215.1050 0.0000 216.6950 0.6300 ;
      RECT 213.1050 0.0000 214.6950 0.6300 ;
      RECT 211.1050 0.0000 212.6950 0.6300 ;
      RECT 209.1050 0.0000 210.6950 0.6300 ;
      RECT 207.1050 0.0000 208.6950 0.6300 ;
      RECT 205.1050 0.0000 206.6950 0.6300 ;
      RECT 203.1050 0.0000 204.6950 0.6300 ;
      RECT 201.1050 0.0000 202.6950 0.6300 ;
      RECT 199.1050 0.0000 200.6950 0.6300 ;
      RECT 197.1050 0.0000 198.6950 0.6300 ;
      RECT 195.1050 0.0000 196.6950 0.6300 ;
      RECT 193.1050 0.0000 194.6950 0.6300 ;
      RECT 191.1050 0.0000 192.6950 0.6300 ;
      RECT 189.1050 0.0000 190.6950 0.6300 ;
      RECT 187.1050 0.0000 188.6950 0.6300 ;
      RECT 185.1050 0.0000 186.6950 0.6300 ;
      RECT 183.1050 0.0000 184.6950 0.6300 ;
      RECT 181.1050 0.0000 182.6950 0.6300 ;
      RECT 179.1050 0.0000 180.6950 0.6300 ;
      RECT 177.1050 0.0000 178.6950 0.6300 ;
      RECT 175.1050 0.0000 176.6950 0.6300 ;
      RECT 173.1050 0.0000 174.6950 0.6300 ;
      RECT 171.1050 0.0000 172.6950 0.6300 ;
      RECT 169.1050 0.0000 170.6950 0.6300 ;
      RECT 167.1050 0.0000 168.6950 0.6300 ;
      RECT 165.1050 0.0000 166.6950 0.6300 ;
      RECT 163.1050 0.0000 164.6950 0.6300 ;
      RECT 161.1050 0.0000 162.6950 0.6300 ;
      RECT 159.1050 0.0000 160.6950 0.6300 ;
      RECT 157.1050 0.0000 158.6950 0.6300 ;
      RECT 155.1050 0.0000 156.6950 0.6300 ;
      RECT 153.1050 0.0000 154.6950 0.6300 ;
      RECT 151.1050 0.0000 152.6950 0.6300 ;
      RECT 149.1050 0.0000 150.6950 0.6300 ;
      RECT 147.1050 0.0000 148.6950 0.6300 ;
      RECT 145.1050 0.0000 146.6950 0.6300 ;
      RECT 143.1050 0.0000 144.6950 0.6300 ;
      RECT 141.1050 0.0000 142.6950 0.6300 ;
      RECT 139.1050 0.0000 140.6950 0.6300 ;
      RECT 137.1050 0.0000 138.6950 0.6300 ;
      RECT 135.1050 0.0000 136.6950 0.6300 ;
      RECT 133.1050 0.0000 134.6950 0.6300 ;
      RECT 131.1050 0.0000 132.6950 0.6300 ;
      RECT 129.1050 0.0000 130.6950 0.6300 ;
      RECT 127.1050 0.0000 128.6950 0.6300 ;
      RECT 125.1050 0.0000 126.6950 0.6300 ;
      RECT 123.1050 0.0000 124.6950 0.6300 ;
      RECT 121.1050 0.0000 122.6950 0.6300 ;
      RECT 119.1050 0.0000 120.6950 0.6300 ;
      RECT 117.1050 0.0000 118.6950 0.6300 ;
      RECT 115.1050 0.0000 116.6950 0.6300 ;
      RECT 113.1050 0.0000 114.6950 0.6300 ;
      RECT 111.1050 0.0000 112.6950 0.6300 ;
      RECT 0.0000 0.0000 110.6950 0.6300 ;
    LAYER M2 ;
      RECT 0.0000 390.0100 540.0000 540.0000 ;
      RECT 0.6800 389.5900 540.0000 390.0100 ;
      RECT 0.0000 387.0100 540.0000 389.5900 ;
      RECT 0.6800 386.5900 540.0000 387.0100 ;
      RECT 0.0000 384.0100 540.0000 386.5900 ;
      RECT 0.6800 383.5900 540.0000 384.0100 ;
      RECT 0.0000 381.0100 540.0000 383.5900 ;
      RECT 0.6800 380.5900 540.0000 381.0100 ;
      RECT 0.0000 378.0100 540.0000 380.5900 ;
      RECT 0.6800 377.5900 540.0000 378.0100 ;
      RECT 0.0000 375.0100 540.0000 377.5900 ;
      RECT 0.6800 374.5900 540.0000 375.0100 ;
      RECT 0.0000 372.0100 540.0000 374.5900 ;
      RECT 0.6800 371.5900 540.0000 372.0100 ;
      RECT 0.0000 369.0100 540.0000 371.5900 ;
      RECT 0.6800 368.5900 540.0000 369.0100 ;
      RECT 0.0000 366.0100 540.0000 368.5900 ;
      RECT 0.6800 365.5900 540.0000 366.0100 ;
      RECT 0.0000 363.0100 540.0000 365.5900 ;
      RECT 0.6800 362.5900 540.0000 363.0100 ;
      RECT 0.0000 360.0100 540.0000 362.5900 ;
      RECT 0.6800 359.5900 540.0000 360.0100 ;
      RECT 0.0000 357.0100 540.0000 359.5900 ;
      RECT 0.6800 356.5900 540.0000 357.0100 ;
      RECT 0.0000 354.0100 540.0000 356.5900 ;
      RECT 0.6800 353.5900 540.0000 354.0100 ;
      RECT 0.0000 351.0100 540.0000 353.5900 ;
      RECT 0.6800 350.5900 540.0000 351.0100 ;
      RECT 0.0000 348.0100 540.0000 350.5900 ;
      RECT 0.6800 347.5900 540.0000 348.0100 ;
      RECT 0.0000 345.0100 540.0000 347.5900 ;
      RECT 0.6800 344.5900 540.0000 345.0100 ;
      RECT 0.0000 342.0100 540.0000 344.5900 ;
      RECT 0.6800 341.5900 540.0000 342.0100 ;
      RECT 0.0000 339.0100 540.0000 341.5900 ;
      RECT 0.6800 338.5900 540.0000 339.0100 ;
      RECT 0.0000 336.0100 540.0000 338.5900 ;
      RECT 0.6800 335.5900 540.0000 336.0100 ;
      RECT 0.0000 333.0100 540.0000 335.5900 ;
      RECT 0.6800 332.5900 540.0000 333.0100 ;
      RECT 0.0000 330.0100 540.0000 332.5900 ;
      RECT 0.6800 329.5900 540.0000 330.0100 ;
      RECT 0.0000 327.0100 540.0000 329.5900 ;
      RECT 0.6800 326.5900 540.0000 327.0100 ;
      RECT 0.0000 324.0100 540.0000 326.5900 ;
      RECT 0.6800 323.5900 540.0000 324.0100 ;
      RECT 0.0000 321.0100 540.0000 323.5900 ;
      RECT 0.6800 320.5900 540.0000 321.0100 ;
      RECT 0.0000 318.0100 540.0000 320.5900 ;
      RECT 0.6800 317.5900 540.0000 318.0100 ;
      RECT 0.0000 315.0100 540.0000 317.5900 ;
      RECT 0.6800 314.5900 540.0000 315.0100 ;
      RECT 0.0000 312.0100 540.0000 314.5900 ;
      RECT 0.6800 311.5900 540.0000 312.0100 ;
      RECT 0.0000 309.0100 540.0000 311.5900 ;
      RECT 0.6800 308.5900 540.0000 309.0100 ;
      RECT 0.0000 306.0100 540.0000 308.5900 ;
      RECT 0.6800 305.5900 540.0000 306.0100 ;
      RECT 0.0000 303.0100 540.0000 305.5900 ;
      RECT 0.6800 302.5900 540.0000 303.0100 ;
      RECT 0.0000 300.0100 540.0000 302.5900 ;
      RECT 0.6800 299.5900 540.0000 300.0100 ;
      RECT 0.0000 297.0100 540.0000 299.5900 ;
      RECT 0.6800 296.5900 540.0000 297.0100 ;
      RECT 0.0000 294.0100 540.0000 296.5900 ;
      RECT 0.6800 293.5900 540.0000 294.0100 ;
      RECT 0.0000 291.0100 540.0000 293.5900 ;
      RECT 0.6800 290.5900 540.0000 291.0100 ;
      RECT 0.0000 288.0100 540.0000 290.5900 ;
      RECT 0.6800 287.5900 540.0000 288.0100 ;
      RECT 0.0000 285.0100 540.0000 287.5900 ;
      RECT 0.6800 284.5900 540.0000 285.0100 ;
      RECT 0.0000 282.0100 540.0000 284.5900 ;
      RECT 0.6800 281.5900 540.0000 282.0100 ;
      RECT 0.0000 279.0100 540.0000 281.5900 ;
      RECT 0.6800 278.5900 540.0000 279.0100 ;
      RECT 0.0000 276.0100 540.0000 278.5900 ;
      RECT 0.6800 275.5900 540.0000 276.0100 ;
      RECT 0.0000 273.0100 540.0000 275.5900 ;
      RECT 0.6800 272.5900 540.0000 273.0100 ;
      RECT 0.0000 270.0100 540.0000 272.5900 ;
      RECT 0.6800 269.5900 540.0000 270.0100 ;
      RECT 0.0000 267.0100 540.0000 269.5900 ;
      RECT 0.6800 266.5900 540.0000 267.0100 ;
      RECT 0.0000 264.0100 540.0000 266.5900 ;
      RECT 0.6800 263.5900 540.0000 264.0100 ;
      RECT 0.0000 261.0100 540.0000 263.5900 ;
      RECT 0.6800 260.5900 540.0000 261.0100 ;
      RECT 0.0000 258.0100 540.0000 260.5900 ;
      RECT 0.6800 257.5900 540.0000 258.0100 ;
      RECT 0.0000 255.0100 540.0000 257.5900 ;
      RECT 0.6800 254.5900 540.0000 255.0100 ;
      RECT 0.0000 252.0100 540.0000 254.5900 ;
      RECT 0.6800 251.5900 540.0000 252.0100 ;
      RECT 0.0000 249.0100 540.0000 251.5900 ;
      RECT 0.6800 248.5900 540.0000 249.0100 ;
      RECT 0.0000 246.0100 540.0000 248.5900 ;
      RECT 0.6800 245.5900 540.0000 246.0100 ;
      RECT 0.0000 243.0100 540.0000 245.5900 ;
      RECT 0.6800 242.5900 540.0000 243.0100 ;
      RECT 0.0000 240.0100 540.0000 242.5900 ;
      RECT 0.6800 239.5900 540.0000 240.0100 ;
      RECT 0.0000 237.0100 540.0000 239.5900 ;
      RECT 0.6800 236.5900 540.0000 237.0100 ;
      RECT 0.0000 234.0100 540.0000 236.5900 ;
      RECT 0.6800 233.5900 540.0000 234.0100 ;
      RECT 0.0000 231.0100 540.0000 233.5900 ;
      RECT 0.6800 230.5900 540.0000 231.0100 ;
      RECT 0.0000 228.0100 540.0000 230.5900 ;
      RECT 0.6800 227.5900 540.0000 228.0100 ;
      RECT 0.0000 225.0100 540.0000 227.5900 ;
      RECT 0.6800 224.5900 540.0000 225.0100 ;
      RECT 0.0000 222.0100 540.0000 224.5900 ;
      RECT 0.6800 221.5900 540.0000 222.0100 ;
      RECT 0.0000 219.0100 540.0000 221.5900 ;
      RECT 0.6800 218.5900 540.0000 219.0100 ;
      RECT 0.0000 216.0100 540.0000 218.5900 ;
      RECT 0.6800 215.5900 540.0000 216.0100 ;
      RECT 0.0000 213.0100 540.0000 215.5900 ;
      RECT 0.6800 212.5900 540.0000 213.0100 ;
      RECT 0.0000 210.0100 540.0000 212.5900 ;
      RECT 0.6800 209.5900 540.0000 210.0100 ;
      RECT 0.0000 207.0100 540.0000 209.5900 ;
      RECT 0.6800 206.5900 540.0000 207.0100 ;
      RECT 0.0000 204.0100 540.0000 206.5900 ;
      RECT 0.6800 203.5900 540.0000 204.0100 ;
      RECT 0.0000 201.0100 540.0000 203.5900 ;
      RECT 0.6800 200.5900 540.0000 201.0100 ;
      RECT 0.0000 198.0100 540.0000 200.5900 ;
      RECT 0.6800 197.5900 540.0000 198.0100 ;
      RECT 0.0000 195.0100 540.0000 197.5900 ;
      RECT 0.6800 194.5900 540.0000 195.0100 ;
      RECT 0.0000 192.0100 540.0000 194.5900 ;
      RECT 0.6800 191.5900 540.0000 192.0100 ;
      RECT 0.0000 189.0100 540.0000 191.5900 ;
      RECT 0.6800 188.5900 540.0000 189.0100 ;
      RECT 0.0000 186.0100 540.0000 188.5900 ;
      RECT 0.6800 185.5900 540.0000 186.0100 ;
      RECT 0.0000 183.0100 540.0000 185.5900 ;
      RECT 0.6800 182.5900 540.0000 183.0100 ;
      RECT 0.0000 180.0100 540.0000 182.5900 ;
      RECT 0.6800 179.5900 540.0000 180.0100 ;
      RECT 0.0000 177.0100 540.0000 179.5900 ;
      RECT 0.6800 176.5900 540.0000 177.0100 ;
      RECT 0.0000 174.0100 540.0000 176.5900 ;
      RECT 0.6800 173.5900 540.0000 174.0100 ;
      RECT 0.0000 171.0100 540.0000 173.5900 ;
      RECT 0.6800 170.5900 540.0000 171.0100 ;
      RECT 0.0000 168.0100 540.0000 170.5900 ;
      RECT 0.6800 167.5900 540.0000 168.0100 ;
      RECT 0.0000 165.0100 540.0000 167.5900 ;
      RECT 0.6800 164.5900 540.0000 165.0100 ;
      RECT 0.0000 162.0100 540.0000 164.5900 ;
      RECT 0.6800 161.5900 540.0000 162.0100 ;
      RECT 0.0000 159.0100 540.0000 161.5900 ;
      RECT 0.6800 158.5900 540.0000 159.0100 ;
      RECT 0.0000 156.0100 540.0000 158.5900 ;
      RECT 0.6800 155.5900 540.0000 156.0100 ;
      RECT 0.0000 153.0100 540.0000 155.5900 ;
      RECT 0.6800 152.5900 540.0000 153.0100 ;
      RECT 0.0000 150.0100 540.0000 152.5900 ;
      RECT 0.6800 149.5900 540.0000 150.0100 ;
      RECT 0.0000 0.0000 540.0000 149.5900 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 540.0000 540.0000 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 540.0000 540.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 540.0000 540.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 540.0000 540.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 540.0000 540.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 540.0000 540.0000 ;
  END
END core

END LIBRARY
