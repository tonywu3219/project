##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 16:56:14 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16_64b
  CLASS BLOCK ;
  SIZE 290.0000 BY 290.0000 ;
  FOREIGN sram_w16_64b 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 152.7500 0.5200 152.8500 ;
    END
  END CLK
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.8500 0.0000 270.9500 0.5200 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 266.8500 0.0000 266.9500 0.5200 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.8500 0.0000 262.9500 0.5200 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.8500 0.0000 258.9500 0.5200 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 254.8500 0.0000 254.9500 0.5200 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.8500 0.0000 250.9500 0.5200 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.8500 0.0000 246.9500 0.5200 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 242.8500 0.0000 242.9500 0.5200 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.8500 0.0000 238.9500 0.5200 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.8500 0.0000 234.9500 0.5200 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.8500 0.0000 230.9500 0.5200 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.8500 0.0000 226.9500 0.5200 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.8500 0.0000 222.9500 0.5200 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.8500 0.0000 218.9500 0.5200 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.8500 0.0000 214.9500 0.5200 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.8500 0.0000 210.9500 0.5200 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.8500 0.0000 206.9500 0.5200 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.8500 0.0000 202.9500 0.5200 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.8500 0.0000 198.9500 0.5200 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.8500 0.0000 194.9500 0.5200 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.8500 0.0000 190.9500 0.5200 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.8500 0.0000 186.9500 0.5200 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.8500 0.0000 182.9500 0.5200 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.8500 0.0000 178.9500 0.5200 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.8500 0.0000 174.9500 0.5200 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.8500 0.0000 170.9500 0.5200 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.8500 0.0000 166.9500 0.5200 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.8500 0.0000 162.9500 0.5200 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.8500 0.0000 158.9500 0.5200 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.8500 0.0000 154.9500 0.5200 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.8500 0.0000 150.9500 0.5200 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.8500 0.0000 146.9500 0.5200 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.8500 0.0000 142.9500 0.5200 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.8500 0.0000 138.9500 0.5200 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.8500 0.0000 134.9500 0.5200 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.8500 0.0000 130.9500 0.5200 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.8500 0.0000 126.9500 0.5200 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.8500 0.0000 122.9500 0.5200 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.8500 0.0000 118.9500 0.5200 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.8500 0.0000 114.9500 0.5200 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.8500 0.0000 110.9500 0.5200 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.8500 0.0000 106.9500 0.5200 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.8500 0.0000 102.9500 0.5200 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.8500 0.0000 98.9500 0.5200 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.8500 0.0000 94.9500 0.5200 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.8500 0.0000 90.9500 0.5200 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.8500 0.0000 86.9500 0.5200 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.8500 0.0000 82.9500 0.5200 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.8500 0.0000 78.9500 0.5200 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.8500 0.0000 74.9500 0.5200 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.8500 0.0000 70.9500 0.5200 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.8500 0.0000 66.9500 0.5200 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.8500 0.0000 62.9500 0.5200 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.8500 0.0000 58.9500 0.5200 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.8500 0.0000 54.9500 0.5200 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.8500 0.0000 50.9500 0.5200 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8500 0.0000 46.9500 0.5200 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.8500 0.0000 42.9500 0.5200 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.8500 0.0000 38.9500 0.5200 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.8500 0.0000 34.9500 0.5200 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.8500 0.0000 30.9500 0.5200 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.8500 0.0000 26.9500 0.5200 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.8500 0.0000 22.9500 0.5200 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.8500 0.0000 18.9500 0.5200 ;
    END
  END D[0]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.8500 289.4800 270.9500 290.0000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 266.8500 289.4800 266.9500 290.0000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.8500 289.4800 262.9500 290.0000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.8500 289.4800 258.9500 290.0000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 254.8500 289.4800 254.9500 290.0000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.8500 289.4800 250.9500 290.0000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.8500 289.4800 246.9500 290.0000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 242.8500 289.4800 242.9500 290.0000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.8500 289.4800 238.9500 290.0000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.8500 289.4800 234.9500 290.0000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.8500 289.4800 230.9500 290.0000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.8500 289.4800 226.9500 290.0000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.8500 289.4800 222.9500 290.0000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.8500 289.4800 218.9500 290.0000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.8500 289.4800 214.9500 290.0000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.8500 289.4800 210.9500 290.0000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.8500 289.4800 206.9500 290.0000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.8500 289.4800 202.9500 290.0000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.8500 289.4800 198.9500 290.0000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.8500 289.4800 194.9500 290.0000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.8500 289.4800 190.9500 290.0000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.8500 289.4800 186.9500 290.0000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.8500 289.4800 182.9500 290.0000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.8500 289.4800 178.9500 290.0000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.8500 289.4800 174.9500 290.0000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.8500 289.4800 170.9500 290.0000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.8500 289.4800 166.9500 290.0000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.8500 289.4800 162.9500 290.0000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.8500 289.4800 158.9500 290.0000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.8500 289.4800 154.9500 290.0000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.8500 289.4800 150.9500 290.0000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.8500 289.4800 146.9500 290.0000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.8500 289.4800 142.9500 290.0000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.8500 289.4800 138.9500 290.0000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.8500 289.4800 134.9500 290.0000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.8500 289.4800 130.9500 290.0000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.8500 289.4800 126.9500 290.0000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.8500 289.4800 122.9500 290.0000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.8500 289.4800 118.9500 290.0000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.8500 289.4800 114.9500 290.0000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.8500 289.4800 110.9500 290.0000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.8500 289.4800 106.9500 290.0000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.8500 289.4800 102.9500 290.0000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.8500 289.4800 98.9500 290.0000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.8500 289.4800 94.9500 290.0000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.8500 289.4800 90.9500 290.0000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.8500 289.4800 86.9500 290.0000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.8500 289.4800 82.9500 290.0000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.8500 289.4800 78.9500 290.0000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.8500 289.4800 74.9500 290.0000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.8500 289.4800 70.9500 290.0000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.8500 289.4800 66.9500 290.0000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.8500 289.4800 62.9500 290.0000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.8500 289.4800 58.9500 290.0000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.8500 289.4800 54.9500 290.0000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.8500 289.4800 50.9500 290.0000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8500 289.4800 46.9500 290.0000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.8500 289.4800 42.9500 290.0000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.8500 289.4800 38.9500 290.0000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.8500 289.4800 34.9500 290.0000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.8500 289.4800 30.9500 290.0000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.8500 289.4800 26.9500 290.0000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.8500 289.4800 22.9500 290.0000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.8500 289.4800 18.9500 290.0000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 148.7500 0.5200 148.8500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 156.7500 0.5200 156.8500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 144.7500 0.5200 144.8500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 140.7500 0.5200 140.8500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 136.7500 0.5200 136.8500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 132.7500 0.5200 132.8500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 35.5450 10.0000 37.5450 280.0000 ;
        RECT 27.0300 10.0000 29.0300 280.0000 ;
        RECT 18.5150 10.0000 20.5150 280.0000 ;
        RECT 10.0000 10.0000 12.0000 280.0000 ;
        RECT 52.5750 10.0000 54.5750 280.0000 ;
        RECT 44.0600 10.0000 46.0600 280.0000 ;
        RECT 61.0900 10.0000 63.0900 280.0000 ;
        RECT 69.6050 10.0000 71.6050 280.0000 ;
        RECT 78.1200 10.0000 80.1200 280.0000 ;
        RECT 86.6350 10.0000 88.6350 280.0000 ;
        RECT 95.1500 10.0000 97.1500 280.0000 ;
        RECT 103.6650 10.0000 105.6650 280.0000 ;
        RECT 112.1800 10.0000 114.1800 280.0000 ;
        RECT 120.6950 10.0000 122.6950 280.0000 ;
        RECT 129.2100 10.0000 131.2100 280.0000 ;
        RECT 137.7250 10.0000 139.7250 280.0000 ;
        RECT 180.3000 10.0000 182.3000 280.0000 ;
        RECT 146.2400 10.0000 148.2400 280.0000 ;
        RECT 154.7550 10.0000 156.7550 280.0000 ;
        RECT 163.2700 10.0000 165.2700 280.0000 ;
        RECT 171.7850 10.0000 173.7850 280.0000 ;
        RECT 188.8150 10.0000 190.8150 280.0000 ;
        RECT 197.3300 10.0000 199.3300 280.0000 ;
        RECT 205.8450 10.0000 207.8450 280.0000 ;
        RECT 214.3600 10.0000 216.3600 280.0000 ;
        RECT 222.8750 10.0000 224.8750 280.0000 ;
        RECT 231.3900 10.0000 233.3900 280.0000 ;
        RECT 239.9050 10.0000 241.9050 280.0000 ;
        RECT 248.4200 10.0000 250.4200 280.0000 ;
        RECT 265.4500 10.0000 267.4500 280.0000 ;
        RECT 256.9350 10.0000 258.9350 280.0000 ;
        RECT 273.9650 10.0000 275.9650 280.0000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 14.0000 10.0000 16.0000 280.0000 ;
        RECT 22.5150 10.0000 24.5150 280.0000 ;
        RECT 31.0300 10.0000 33.0300 280.0000 ;
        RECT 48.0600 10.0000 50.0600 280.0000 ;
        RECT 39.5450 10.0000 41.5450 280.0000 ;
        RECT 65.0900 10.0000 67.0900 280.0000 ;
        RECT 56.5750 10.0000 58.5750 280.0000 ;
        RECT 107.6650 10.0000 109.6650 280.0000 ;
        RECT 82.1200 10.0000 84.1200 280.0000 ;
        RECT 73.6050 10.0000 75.6050 280.0000 ;
        RECT 99.1500 10.0000 101.1500 280.0000 ;
        RECT 90.6350 10.0000 92.6350 280.0000 ;
        RECT 124.6950 10.0000 126.6950 280.0000 ;
        RECT 116.1800 10.0000 118.1800 280.0000 ;
        RECT 133.2100 10.0000 135.2100 280.0000 ;
        RECT 141.7250 10.0000 143.7250 280.0000 ;
        RECT 158.7550 10.0000 160.7550 280.0000 ;
        RECT 150.2400 10.0000 152.2400 280.0000 ;
        RECT 175.7850 10.0000 177.7850 280.0000 ;
        RECT 167.2700 10.0000 169.2700 280.0000 ;
        RECT 192.8150 10.0000 194.8150 280.0000 ;
        RECT 184.3000 10.0000 186.3000 280.0000 ;
        RECT 209.8450 10.0000 211.8450 280.0000 ;
        RECT 201.3300 10.0000 203.3300 280.0000 ;
        RECT 252.4200 10.0000 254.4200 280.0000 ;
        RECT 235.3900 10.0000 237.3900 280.0000 ;
        RECT 226.8750 10.0000 228.8750 280.0000 ;
        RECT 218.3600 10.0000 220.3600 280.0000 ;
        RECT 243.9050 10.0000 245.9050 280.0000 ;
        RECT 277.9650 10.0000 279.9650 280.0000 ;
        RECT 269.4500 10.0000 271.4500 280.0000 ;
        RECT 260.9350 10.0000 262.9350 280.0000 ;
        RECT 14.0000 9.8350 16.0000 10.1650 ;
        RECT 22.5150 9.8350 24.5150 10.1650 ;
        RECT 31.0300 9.8350 33.0300 10.1650 ;
        RECT 39.5450 9.8350 41.5450 10.1650 ;
        RECT 48.0600 9.8350 50.0600 10.1650 ;
        RECT 56.5750 9.8350 58.5750 10.1650 ;
        RECT 65.0900 9.8350 67.0900 10.1650 ;
        RECT 107.6650 9.8350 109.6650 10.1650 ;
        RECT 73.6050 9.8350 75.6050 10.1650 ;
        RECT 82.1200 9.8350 84.1200 10.1650 ;
        RECT 99.1500 9.8350 101.1500 10.1650 ;
        RECT 90.6350 9.8350 92.6350 10.1650 ;
        RECT 116.1800 9.8350 118.1800 10.1650 ;
        RECT 124.6950 9.8350 126.6950 10.1650 ;
        RECT 133.2100 9.8350 135.2100 10.1650 ;
        RECT 141.7250 9.8350 143.7250 10.1650 ;
        RECT 150.2400 9.8350 152.2400 10.1650 ;
        RECT 158.7550 9.8350 160.7550 10.1650 ;
        RECT 167.2700 9.8350 169.2700 10.1650 ;
        RECT 175.7850 9.8350 177.7850 10.1650 ;
        RECT 184.3000 9.8350 186.3000 10.1650 ;
        RECT 192.8150 9.8350 194.8150 10.1650 ;
        RECT 201.3300 9.8350 203.3300 10.1650 ;
        RECT 209.8450 9.8350 211.8450 10.1650 ;
        RECT 252.4200 9.8350 254.4200 10.1650 ;
        RECT 235.3900 9.8350 237.3900 10.1650 ;
        RECT 218.3600 9.8350 220.3600 10.1650 ;
        RECT 226.8750 9.8350 228.8750 10.1650 ;
        RECT 243.9050 9.8350 245.9050 10.1650 ;
        RECT 260.9350 9.8350 262.9350 10.1650 ;
        RECT 269.4500 9.8350 271.4500 10.1650 ;
        RECT 277.9650 9.8350 279.9650 10.1650 ;
        RECT 14.0000 279.8350 16.0000 280.1650 ;
        RECT 22.5150 279.8350 24.5150 280.1650 ;
        RECT 31.0300 279.8350 33.0300 280.1650 ;
        RECT 39.5450 279.8350 41.5450 280.1650 ;
        RECT 48.0600 279.8350 50.0600 280.1650 ;
        RECT 56.5750 279.8350 58.5750 280.1650 ;
        RECT 65.0900 279.8350 67.0900 280.1650 ;
        RECT 107.6650 279.8350 109.6650 280.1650 ;
        RECT 73.6050 279.8350 75.6050 280.1650 ;
        RECT 82.1200 279.8350 84.1200 280.1650 ;
        RECT 99.1500 279.8350 101.1500 280.1650 ;
        RECT 90.6350 279.8350 92.6350 280.1650 ;
        RECT 116.1800 279.8350 118.1800 280.1650 ;
        RECT 124.6950 279.8350 126.6950 280.1650 ;
        RECT 133.2100 279.8350 135.2100 280.1650 ;
        RECT 141.7250 279.8350 143.7250 280.1650 ;
        RECT 150.2400 279.8350 152.2400 280.1650 ;
        RECT 158.7550 279.8350 160.7550 280.1650 ;
        RECT 167.2700 279.8350 169.2700 280.1650 ;
        RECT 175.7850 279.8350 177.7850 280.1650 ;
        RECT 184.3000 279.8350 186.3000 280.1650 ;
        RECT 192.8150 279.8350 194.8150 280.1650 ;
        RECT 201.3300 279.8350 203.3300 280.1650 ;
        RECT 209.8450 279.8350 211.8450 280.1650 ;
        RECT 252.4200 279.8350 254.4200 280.1650 ;
        RECT 235.3900 279.8350 237.3900 280.1650 ;
        RECT 218.3600 279.8350 220.3600 280.1650 ;
        RECT 226.8750 279.8350 228.8750 280.1650 ;
        RECT 243.9050 279.8350 245.9050 280.1650 ;
        RECT 260.9350 279.8350 262.9350 280.1650 ;
        RECT 269.4500 279.8350 271.4500 280.1650 ;
        RECT 277.9650 279.8350 279.9650 280.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 290.0000 290.0000 ;
    LAYER M2 ;
      RECT 271.0500 289.3800 290.0000 290.0000 ;
      RECT 267.0500 289.3800 270.7500 290.0000 ;
      RECT 263.0500 289.3800 266.7500 290.0000 ;
      RECT 259.0500 289.3800 262.7500 290.0000 ;
      RECT 255.0500 289.3800 258.7500 290.0000 ;
      RECT 251.0500 289.3800 254.7500 290.0000 ;
      RECT 247.0500 289.3800 250.7500 290.0000 ;
      RECT 243.0500 289.3800 246.7500 290.0000 ;
      RECT 239.0500 289.3800 242.7500 290.0000 ;
      RECT 235.0500 289.3800 238.7500 290.0000 ;
      RECT 231.0500 289.3800 234.7500 290.0000 ;
      RECT 227.0500 289.3800 230.7500 290.0000 ;
      RECT 223.0500 289.3800 226.7500 290.0000 ;
      RECT 219.0500 289.3800 222.7500 290.0000 ;
      RECT 215.0500 289.3800 218.7500 290.0000 ;
      RECT 211.0500 289.3800 214.7500 290.0000 ;
      RECT 207.0500 289.3800 210.7500 290.0000 ;
      RECT 203.0500 289.3800 206.7500 290.0000 ;
      RECT 199.0500 289.3800 202.7500 290.0000 ;
      RECT 195.0500 289.3800 198.7500 290.0000 ;
      RECT 191.0500 289.3800 194.7500 290.0000 ;
      RECT 187.0500 289.3800 190.7500 290.0000 ;
      RECT 183.0500 289.3800 186.7500 290.0000 ;
      RECT 179.0500 289.3800 182.7500 290.0000 ;
      RECT 175.0500 289.3800 178.7500 290.0000 ;
      RECT 171.0500 289.3800 174.7500 290.0000 ;
      RECT 167.0500 289.3800 170.7500 290.0000 ;
      RECT 163.0500 289.3800 166.7500 290.0000 ;
      RECT 159.0500 289.3800 162.7500 290.0000 ;
      RECT 155.0500 289.3800 158.7500 290.0000 ;
      RECT 151.0500 289.3800 154.7500 290.0000 ;
      RECT 147.0500 289.3800 150.7500 290.0000 ;
      RECT 143.0500 289.3800 146.7500 290.0000 ;
      RECT 139.0500 289.3800 142.7500 290.0000 ;
      RECT 135.0500 289.3800 138.7500 290.0000 ;
      RECT 131.0500 289.3800 134.7500 290.0000 ;
      RECT 127.0500 289.3800 130.7500 290.0000 ;
      RECT 123.0500 289.3800 126.7500 290.0000 ;
      RECT 119.0500 289.3800 122.7500 290.0000 ;
      RECT 115.0500 289.3800 118.7500 290.0000 ;
      RECT 111.0500 289.3800 114.7500 290.0000 ;
      RECT 107.0500 289.3800 110.7500 290.0000 ;
      RECT 103.0500 289.3800 106.7500 290.0000 ;
      RECT 99.0500 289.3800 102.7500 290.0000 ;
      RECT 95.0500 289.3800 98.7500 290.0000 ;
      RECT 91.0500 289.3800 94.7500 290.0000 ;
      RECT 87.0500 289.3800 90.7500 290.0000 ;
      RECT 83.0500 289.3800 86.7500 290.0000 ;
      RECT 79.0500 289.3800 82.7500 290.0000 ;
      RECT 75.0500 289.3800 78.7500 290.0000 ;
      RECT 71.0500 289.3800 74.7500 290.0000 ;
      RECT 67.0500 289.3800 70.7500 290.0000 ;
      RECT 63.0500 289.3800 66.7500 290.0000 ;
      RECT 59.0500 289.3800 62.7500 290.0000 ;
      RECT 55.0500 289.3800 58.7500 290.0000 ;
      RECT 51.0500 289.3800 54.7500 290.0000 ;
      RECT 47.0500 289.3800 50.7500 290.0000 ;
      RECT 43.0500 289.3800 46.7500 290.0000 ;
      RECT 39.0500 289.3800 42.7500 290.0000 ;
      RECT 35.0500 289.3800 38.7500 290.0000 ;
      RECT 31.0500 289.3800 34.7500 290.0000 ;
      RECT 27.0500 289.3800 30.7500 290.0000 ;
      RECT 23.0500 289.3800 26.7500 290.0000 ;
      RECT 19.0500 289.3800 22.7500 290.0000 ;
      RECT 0.0000 289.3800 18.7500 290.0000 ;
      RECT 0.0000 0.6200 290.0000 289.3800 ;
      RECT 271.0500 0.0000 290.0000 0.6200 ;
      RECT 267.0500 0.0000 270.7500 0.6200 ;
      RECT 263.0500 0.0000 266.7500 0.6200 ;
      RECT 259.0500 0.0000 262.7500 0.6200 ;
      RECT 255.0500 0.0000 258.7500 0.6200 ;
      RECT 251.0500 0.0000 254.7500 0.6200 ;
      RECT 247.0500 0.0000 250.7500 0.6200 ;
      RECT 243.0500 0.0000 246.7500 0.6200 ;
      RECT 239.0500 0.0000 242.7500 0.6200 ;
      RECT 235.0500 0.0000 238.7500 0.6200 ;
      RECT 231.0500 0.0000 234.7500 0.6200 ;
      RECT 227.0500 0.0000 230.7500 0.6200 ;
      RECT 223.0500 0.0000 226.7500 0.6200 ;
      RECT 219.0500 0.0000 222.7500 0.6200 ;
      RECT 215.0500 0.0000 218.7500 0.6200 ;
      RECT 211.0500 0.0000 214.7500 0.6200 ;
      RECT 207.0500 0.0000 210.7500 0.6200 ;
      RECT 203.0500 0.0000 206.7500 0.6200 ;
      RECT 199.0500 0.0000 202.7500 0.6200 ;
      RECT 195.0500 0.0000 198.7500 0.6200 ;
      RECT 191.0500 0.0000 194.7500 0.6200 ;
      RECT 187.0500 0.0000 190.7500 0.6200 ;
      RECT 183.0500 0.0000 186.7500 0.6200 ;
      RECT 179.0500 0.0000 182.7500 0.6200 ;
      RECT 175.0500 0.0000 178.7500 0.6200 ;
      RECT 171.0500 0.0000 174.7500 0.6200 ;
      RECT 167.0500 0.0000 170.7500 0.6200 ;
      RECT 163.0500 0.0000 166.7500 0.6200 ;
      RECT 159.0500 0.0000 162.7500 0.6200 ;
      RECT 155.0500 0.0000 158.7500 0.6200 ;
      RECT 151.0500 0.0000 154.7500 0.6200 ;
      RECT 147.0500 0.0000 150.7500 0.6200 ;
      RECT 143.0500 0.0000 146.7500 0.6200 ;
      RECT 139.0500 0.0000 142.7500 0.6200 ;
      RECT 135.0500 0.0000 138.7500 0.6200 ;
      RECT 131.0500 0.0000 134.7500 0.6200 ;
      RECT 127.0500 0.0000 130.7500 0.6200 ;
      RECT 123.0500 0.0000 126.7500 0.6200 ;
      RECT 119.0500 0.0000 122.7500 0.6200 ;
      RECT 115.0500 0.0000 118.7500 0.6200 ;
      RECT 111.0500 0.0000 114.7500 0.6200 ;
      RECT 107.0500 0.0000 110.7500 0.6200 ;
      RECT 103.0500 0.0000 106.7500 0.6200 ;
      RECT 99.0500 0.0000 102.7500 0.6200 ;
      RECT 95.0500 0.0000 98.7500 0.6200 ;
      RECT 91.0500 0.0000 94.7500 0.6200 ;
      RECT 87.0500 0.0000 90.7500 0.6200 ;
      RECT 83.0500 0.0000 86.7500 0.6200 ;
      RECT 79.0500 0.0000 82.7500 0.6200 ;
      RECT 75.0500 0.0000 78.7500 0.6200 ;
      RECT 71.0500 0.0000 74.7500 0.6200 ;
      RECT 67.0500 0.0000 70.7500 0.6200 ;
      RECT 63.0500 0.0000 66.7500 0.6200 ;
      RECT 59.0500 0.0000 62.7500 0.6200 ;
      RECT 55.0500 0.0000 58.7500 0.6200 ;
      RECT 51.0500 0.0000 54.7500 0.6200 ;
      RECT 47.0500 0.0000 50.7500 0.6200 ;
      RECT 43.0500 0.0000 46.7500 0.6200 ;
      RECT 39.0500 0.0000 42.7500 0.6200 ;
      RECT 35.0500 0.0000 38.7500 0.6200 ;
      RECT 31.0500 0.0000 34.7500 0.6200 ;
      RECT 27.0500 0.0000 30.7500 0.6200 ;
      RECT 23.0500 0.0000 26.7500 0.6200 ;
      RECT 19.0500 0.0000 22.7500 0.6200 ;
      RECT 0.0000 0.0000 18.7500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 156.9500 290.0000 290.0000 ;
      RECT 0.6200 156.6500 290.0000 156.9500 ;
      RECT 0.0000 152.9500 290.0000 156.6500 ;
      RECT 0.6200 152.6500 290.0000 152.9500 ;
      RECT 0.0000 148.9500 290.0000 152.6500 ;
      RECT 0.6200 148.6500 290.0000 148.9500 ;
      RECT 0.0000 144.9500 290.0000 148.6500 ;
      RECT 0.6200 144.6500 290.0000 144.9500 ;
      RECT 0.0000 140.9500 290.0000 144.6500 ;
      RECT 0.6200 140.6500 290.0000 140.9500 ;
      RECT 0.0000 136.9500 290.0000 140.6500 ;
      RECT 0.6200 136.6500 290.0000 136.9500 ;
      RECT 0.0000 132.9500 290.0000 136.6500 ;
      RECT 0.6200 132.6500 290.0000 132.9500 ;
      RECT 0.0000 0.0000 290.0000 132.6500 ;
    LAYER M4 ;
      RECT 0.0000 280.6650 290.0000 290.0000 ;
      RECT 271.9500 280.5000 277.4650 280.6650 ;
      RECT 263.4350 280.5000 268.9500 280.6650 ;
      RECT 254.9200 280.5000 260.4350 280.6650 ;
      RECT 246.4050 280.5000 251.9200 280.6650 ;
      RECT 237.8900 280.5000 243.4050 280.6650 ;
      RECT 229.3750 280.5000 234.8900 280.6650 ;
      RECT 220.8600 280.5000 226.3750 280.6650 ;
      RECT 212.3450 280.5000 217.8600 280.6650 ;
      RECT 203.8300 280.5000 209.3450 280.6650 ;
      RECT 195.3150 280.5000 200.8300 280.6650 ;
      RECT 186.8000 280.5000 192.3150 280.6650 ;
      RECT 178.2850 280.5000 183.8000 280.6650 ;
      RECT 169.7700 280.5000 175.2850 280.6650 ;
      RECT 161.2550 280.5000 166.7700 280.6650 ;
      RECT 152.7400 280.5000 158.2550 280.6650 ;
      RECT 144.2250 280.5000 149.7400 280.6650 ;
      RECT 135.7100 280.5000 141.2250 280.6650 ;
      RECT 127.1950 280.5000 132.7100 280.6650 ;
      RECT 118.6800 280.5000 124.1950 280.6650 ;
      RECT 110.1650 280.5000 115.6800 280.6650 ;
      RECT 101.6500 280.5000 107.1650 280.6650 ;
      RECT 93.1350 280.5000 98.6500 280.6650 ;
      RECT 84.6200 280.5000 90.1350 280.6650 ;
      RECT 76.1050 280.5000 81.6200 280.6650 ;
      RECT 67.5900 280.5000 73.1050 280.6650 ;
      RECT 59.0750 280.5000 64.5900 280.6650 ;
      RECT 50.5600 280.5000 56.0750 280.6650 ;
      RECT 42.0450 280.5000 47.5600 280.6650 ;
      RECT 33.5300 280.5000 39.0450 280.6650 ;
      RECT 25.0150 280.5000 30.5300 280.6650 ;
      RECT 16.5000 280.5000 22.0150 280.6650 ;
      RECT 0.0000 280.5000 13.5000 280.6650 ;
      RECT 276.4650 9.5000 277.4650 280.5000 ;
      RECT 271.9500 9.5000 273.4650 280.5000 ;
      RECT 267.9500 9.5000 268.9500 280.5000 ;
      RECT 263.4350 9.5000 264.9500 280.5000 ;
      RECT 259.4350 9.5000 260.4350 280.5000 ;
      RECT 254.9200 9.5000 256.4350 280.5000 ;
      RECT 250.9200 9.5000 251.9200 280.5000 ;
      RECT 246.4050 9.5000 247.9200 280.5000 ;
      RECT 242.4050 9.5000 243.4050 280.5000 ;
      RECT 237.8900 9.5000 239.4050 280.5000 ;
      RECT 233.8900 9.5000 234.8900 280.5000 ;
      RECT 229.3750 9.5000 230.8900 280.5000 ;
      RECT 225.3750 9.5000 226.3750 280.5000 ;
      RECT 220.8600 9.5000 222.3750 280.5000 ;
      RECT 216.8600 9.5000 217.8600 280.5000 ;
      RECT 212.3450 9.5000 213.8600 280.5000 ;
      RECT 208.3450 9.5000 209.3450 280.5000 ;
      RECT 203.8300 9.5000 205.3450 280.5000 ;
      RECT 199.8300 9.5000 200.8300 280.5000 ;
      RECT 195.3150 9.5000 196.8300 280.5000 ;
      RECT 191.3150 9.5000 192.3150 280.5000 ;
      RECT 186.8000 9.5000 188.3150 280.5000 ;
      RECT 182.8000 9.5000 183.8000 280.5000 ;
      RECT 178.2850 9.5000 179.8000 280.5000 ;
      RECT 174.2850 9.5000 175.2850 280.5000 ;
      RECT 169.7700 9.5000 171.2850 280.5000 ;
      RECT 165.7700 9.5000 166.7700 280.5000 ;
      RECT 161.2550 9.5000 162.7700 280.5000 ;
      RECT 157.2550 9.5000 158.2550 280.5000 ;
      RECT 152.7400 9.5000 154.2550 280.5000 ;
      RECT 148.7400 9.5000 149.7400 280.5000 ;
      RECT 144.2250 9.5000 145.7400 280.5000 ;
      RECT 140.2250 9.5000 141.2250 280.5000 ;
      RECT 135.7100 9.5000 137.2250 280.5000 ;
      RECT 131.7100 9.5000 132.7100 280.5000 ;
      RECT 127.1950 9.5000 128.7100 280.5000 ;
      RECT 123.1950 9.5000 124.1950 280.5000 ;
      RECT 118.6800 9.5000 120.1950 280.5000 ;
      RECT 114.6800 9.5000 115.6800 280.5000 ;
      RECT 110.1650 9.5000 111.6800 280.5000 ;
      RECT 106.1650 9.5000 107.1650 280.5000 ;
      RECT 101.6500 9.5000 103.1650 280.5000 ;
      RECT 97.6500 9.5000 98.6500 280.5000 ;
      RECT 93.1350 9.5000 94.6500 280.5000 ;
      RECT 89.1350 9.5000 90.1350 280.5000 ;
      RECT 84.6200 9.5000 86.1350 280.5000 ;
      RECT 80.6200 9.5000 81.6200 280.5000 ;
      RECT 76.1050 9.5000 77.6200 280.5000 ;
      RECT 72.1050 9.5000 73.1050 280.5000 ;
      RECT 67.5900 9.5000 69.1050 280.5000 ;
      RECT 63.5900 9.5000 64.5900 280.5000 ;
      RECT 59.0750 9.5000 60.5900 280.5000 ;
      RECT 55.0750 9.5000 56.0750 280.5000 ;
      RECT 50.5600 9.5000 52.0750 280.5000 ;
      RECT 46.5600 9.5000 47.5600 280.5000 ;
      RECT 42.0450 9.5000 43.5600 280.5000 ;
      RECT 38.0450 9.5000 39.0450 280.5000 ;
      RECT 33.5300 9.5000 35.0450 280.5000 ;
      RECT 29.5300 9.5000 30.5300 280.5000 ;
      RECT 25.0150 9.5000 26.5300 280.5000 ;
      RECT 21.0150 9.5000 22.0150 280.5000 ;
      RECT 16.5000 9.5000 18.0150 280.5000 ;
      RECT 12.5000 9.5000 13.5000 280.5000 ;
      RECT 0.0000 9.5000 9.5000 280.5000 ;
      RECT 280.4650 9.3350 290.0000 280.6650 ;
      RECT 271.9500 9.3350 277.4650 9.5000 ;
      RECT 263.4350 9.3350 268.9500 9.5000 ;
      RECT 254.9200 9.3350 260.4350 9.5000 ;
      RECT 246.4050 9.3350 251.9200 9.5000 ;
      RECT 237.8900 9.3350 243.4050 9.5000 ;
      RECT 229.3750 9.3350 234.8900 9.5000 ;
      RECT 220.8600 9.3350 226.3750 9.5000 ;
      RECT 212.3450 9.3350 217.8600 9.5000 ;
      RECT 203.8300 9.3350 209.3450 9.5000 ;
      RECT 195.3150 9.3350 200.8300 9.5000 ;
      RECT 186.8000 9.3350 192.3150 9.5000 ;
      RECT 178.2850 9.3350 183.8000 9.5000 ;
      RECT 169.7700 9.3350 175.2850 9.5000 ;
      RECT 161.2550 9.3350 166.7700 9.5000 ;
      RECT 152.7400 9.3350 158.2550 9.5000 ;
      RECT 144.2250 9.3350 149.7400 9.5000 ;
      RECT 135.7100 9.3350 141.2250 9.5000 ;
      RECT 127.1950 9.3350 132.7100 9.5000 ;
      RECT 118.6800 9.3350 124.1950 9.5000 ;
      RECT 110.1650 9.3350 115.6800 9.5000 ;
      RECT 101.6500 9.3350 107.1650 9.5000 ;
      RECT 93.1350 9.3350 98.6500 9.5000 ;
      RECT 84.6200 9.3350 90.1350 9.5000 ;
      RECT 76.1050 9.3350 81.6200 9.5000 ;
      RECT 67.5900 9.3350 73.1050 9.5000 ;
      RECT 59.0750 9.3350 64.5900 9.5000 ;
      RECT 50.5600 9.3350 56.0750 9.5000 ;
      RECT 42.0450 9.3350 47.5600 9.5000 ;
      RECT 33.5300 9.3350 39.0450 9.5000 ;
      RECT 25.0150 9.3350 30.5300 9.5000 ;
      RECT 16.5000 9.3350 22.0150 9.5000 ;
      RECT 0.0000 9.3350 13.5000 9.5000 ;
      RECT 0.0000 0.0000 290.0000 9.3350 ;
  END
END sram_w16_64b

END LIBRARY
