##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar  8 14:33:49 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 570.0000 BY 570.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 282.2550 569.5300 282.3450 570.0000 ;
    END
  END clk
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 559.2550 0.0000 559.3450 0.4700 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 556.2550 0.0000 556.3450 0.4700 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 553.2550 0.0000 553.3450 0.4700 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 550.2550 0.0000 550.3450 0.4700 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 547.2550 0.0000 547.3450 0.4700 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 544.2550 0.0000 544.3450 0.4700 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 541.2550 0.0000 541.3450 0.4700 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 538.2550 0.0000 538.3450 0.4700 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 535.2550 0.0000 535.3450 0.4700 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 532.2550 0.0000 532.3450 0.4700 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 529.2550 0.0000 529.3450 0.4700 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 526.2550 0.0000 526.3450 0.4700 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 523.2550 0.0000 523.3450 0.4700 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 520.2550 0.0000 520.3450 0.4700 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 517.2550 0.0000 517.3450 0.4700 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 514.2550 0.0000 514.3450 0.4700 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 511.2550 0.0000 511.3450 0.4700 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 508.2550 0.0000 508.3450 0.4700 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 505.2550 0.0000 505.3450 0.4700 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 502.2550 0.0000 502.3450 0.4700 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 499.2550 0.0000 499.3450 0.4700 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 496.2550 0.0000 496.3450 0.4700 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 493.2550 0.0000 493.3450 0.4700 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 490.2550 0.0000 490.3450 0.4700 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 484.7500 0.5200 484.8500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 479.7500 0.5200 479.8500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 474.7500 0.5200 474.8500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 469.7500 0.5200 469.8500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 464.7500 0.5200 464.8500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 459.7500 0.5200 459.8500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 454.7500 0.5200 454.8500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 449.7500 0.5200 449.8500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 444.7500 0.5200 444.8500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 439.7500 0.5200 439.8500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 434.7500 0.5200 434.8500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 429.7500 0.5200 429.8500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 424.7500 0.5200 424.8500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 419.7500 0.5200 419.8500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 414.7500 0.5200 414.8500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 409.7500 0.5200 409.8500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 404.7500 0.5200 404.8500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 399.7500 0.5200 399.8500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 394.7500 0.5200 394.8500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 389.7500 0.5200 389.8500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 384.7500 0.5200 384.8500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 379.7500 0.5200 379.8500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 374.7500 0.5200 374.8500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 369.7500 0.5200 369.8500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 364.7500 0.5200 364.8500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 359.7500 0.5200 359.8500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 354.7500 0.5200 354.8500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 349.7500 0.5200 349.8500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 344.7500 0.5200 344.8500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 339.7500 0.5200 339.8500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 334.7500 0.5200 334.8500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 329.7500 0.5200 329.8500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 324.7500 0.5200 324.8500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 319.7500 0.5200 319.8500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 314.7500 0.5200 314.8500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 309.7500 0.5200 309.8500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 304.7500 0.5200 304.8500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 299.7500 0.5200 299.8500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 294.7500 0.5200 294.8500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 289.7500 0.5200 289.8500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 284.7500 0.5200 284.8500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 279.7500 0.5200 279.8500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 274.7500 0.5200 274.8500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 269.7500 0.5200 269.8500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 264.7500 0.5200 264.8500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 259.7500 0.5200 259.8500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 254.7500 0.5200 254.8500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 249.7500 0.5200 249.8500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 244.7500 0.5200 244.8500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 239.7500 0.5200 239.8500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 234.7500 0.5200 234.8500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 229.7500 0.5200 229.8500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 224.7500 0.5200 224.8500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 219.7500 0.5200 219.8500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 214.7500 0.5200 214.8500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 209.7500 0.5200 209.8500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 204.7500 0.5200 204.8500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 199.7500 0.5200 199.8500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 194.7500 0.5200 194.8500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 189.7500 0.5200 189.8500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 184.7500 0.5200 184.8500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 179.7500 0.5200 179.8500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 174.7500 0.5200 174.8500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 169.7500 0.5200 169.8500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 487.2550 0.0000 487.3450 0.4700 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 484.2550 0.0000 484.3450 0.4700 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 481.2550 0.0000 481.3450 0.4700 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 478.2550 0.0000 478.3450 0.4700 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 475.2550 0.0000 475.3450 0.4700 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 472.2550 0.0000 472.3450 0.4700 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 469.2550 0.0000 469.3450 0.4700 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 466.2550 0.0000 466.3450 0.4700 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 463.2550 0.0000 463.3450 0.4700 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 460.2550 0.0000 460.3450 0.4700 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 457.2550 0.0000 457.3450 0.4700 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 454.2550 0.0000 454.3450 0.4700 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 451.2550 0.0000 451.3450 0.4700 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 448.2550 0.0000 448.3450 0.4700 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 445.2550 0.0000 445.3450 0.4700 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 442.2550 0.0000 442.3450 0.4700 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 439.2550 0.0000 439.3450 0.4700 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 436.2550 0.0000 436.3450 0.4700 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 433.2550 0.0000 433.3450 0.4700 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 430.2550 0.0000 430.3450 0.4700 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 427.2550 0.0000 427.3450 0.4700 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 424.2550 0.0000 424.3450 0.4700 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 421.2550 0.0000 421.3450 0.4700 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 418.2550 0.0000 418.3450 0.4700 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 415.2550 0.0000 415.3450 0.4700 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 412.2550 0.0000 412.3450 0.4700 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 409.2550 0.0000 409.3450 0.4700 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 406.2550 0.0000 406.3450 0.4700 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 403.2550 0.0000 403.3450 0.4700 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 400.2550 0.0000 400.3450 0.4700 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 397.2550 0.0000 397.3450 0.4700 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 394.2550 0.0000 394.3450 0.4700 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 391.2550 0.0000 391.3450 0.4700 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 388.2550 0.0000 388.3450 0.4700 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 385.2550 0.0000 385.3450 0.4700 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 382.2550 0.0000 382.3450 0.4700 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 379.2550 0.0000 379.3450 0.4700 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 376.2550 0.0000 376.3450 0.4700 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 373.2550 0.0000 373.3450 0.4700 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 370.2550 0.0000 370.3450 0.4700 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 367.2550 0.0000 367.3450 0.4700 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 364.2550 0.0000 364.3450 0.4700 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 361.2550 0.0000 361.3450 0.4700 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 358.2550 0.0000 358.3450 0.4700 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 355.2550 0.0000 355.3450 0.4700 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 352.2550 0.0000 352.3450 0.4700 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 349.2550 0.0000 349.3450 0.4700 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 346.2550 0.0000 346.3450 0.4700 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 343.2550 0.0000 343.3450 0.4700 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 340.2550 0.0000 340.3450 0.4700 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 337.2550 0.0000 337.3450 0.4700 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 334.2550 0.0000 334.3450 0.4700 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 331.2550 0.0000 331.3450 0.4700 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 328.2550 0.0000 328.3450 0.4700 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 325.2550 0.0000 325.3450 0.4700 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 322.2550 0.0000 322.3450 0.4700 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 319.2550 0.0000 319.3450 0.4700 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 316.2550 0.0000 316.3450 0.4700 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 313.2550 0.0000 313.3450 0.4700 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 310.2550 0.0000 310.3450 0.4700 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 307.2550 0.0000 307.3450 0.4700 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 304.2550 0.0000 304.3450 0.4700 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 301.2550 0.0000 301.3450 0.4700 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 298.2550 0.0000 298.3450 0.4700 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 295.2550 0.0000 295.3450 0.4700 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 292.2550 0.0000 292.3450 0.4700 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 289.2550 0.0000 289.3450 0.4700 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 286.2550 0.0000 286.3450 0.4700 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 283.2550 0.0000 283.3450 0.4700 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 280.2550 0.0000 280.3450 0.4700 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 277.2550 0.0000 277.3450 0.4700 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 274.2550 0.0000 274.3450 0.4700 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 271.2550 0.0000 271.3450 0.4700 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 268.2550 0.0000 268.3450 0.4700 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 265.2550 0.0000 265.3450 0.4700 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 262.2550 0.0000 262.3450 0.4700 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 259.2550 0.0000 259.3450 0.4700 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 256.2550 0.0000 256.3450 0.4700 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 253.2550 0.0000 253.3450 0.4700 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 250.2550 0.0000 250.3450 0.4700 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 247.2550 0.0000 247.3450 0.4700 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 244.2550 0.0000 244.3450 0.4700 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 241.2550 0.0000 241.3450 0.4700 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 238.2550 0.0000 238.3450 0.4700 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 235.2550 0.0000 235.3450 0.4700 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 232.2550 0.0000 232.3450 0.4700 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 229.2550 0.0000 229.3450 0.4700 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 226.2550 0.0000 226.3450 0.4700 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 223.2550 0.0000 223.3450 0.4700 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 220.2550 0.0000 220.3450 0.4700 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 217.2550 0.0000 217.3450 0.4700 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 214.2550 0.0000 214.3450 0.4700 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 211.2550 0.0000 211.3450 0.4700 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 208.2550 0.0000 208.3450 0.4700 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 205.2550 0.0000 205.3450 0.4700 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 202.2550 0.0000 202.3450 0.4700 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 199.2550 0.0000 199.3450 0.4700 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 196.2550 0.0000 196.3450 0.4700 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 193.2550 0.0000 193.3450 0.4700 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 190.2550 0.0000 190.3450 0.4700 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 187.2550 0.0000 187.3450 0.4700 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 184.2550 0.0000 184.3450 0.4700 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 181.2550 0.0000 181.3450 0.4700 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 178.2550 0.0000 178.3450 0.4700 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 175.2550 0.0000 175.3450 0.4700 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 172.2550 0.0000 172.3450 0.4700 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 169.2550 0.0000 169.3450 0.4700 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 166.2550 0.0000 166.3450 0.4700 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 163.2550 0.0000 163.3450 0.4700 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 160.2550 0.0000 160.3450 0.4700 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 157.2550 0.0000 157.3450 0.4700 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 154.2550 0.0000 154.3450 0.4700 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 151.2550 0.0000 151.3450 0.4700 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 148.2550 0.0000 148.3450 0.4700 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 145.2550 0.0000 145.3450 0.4700 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 142.2550 0.0000 142.3450 0.4700 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 139.2550 0.0000 139.3450 0.4700 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 136.2550 0.0000 136.3450 0.4700 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 133.2550 0.0000 133.3450 0.4700 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 130.2550 0.0000 130.3450 0.4700 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 127.2550 0.0000 127.3450 0.4700 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 124.2550 0.0000 124.3450 0.4700 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 121.2550 0.0000 121.3450 0.4700 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 118.2550 0.0000 118.3450 0.4700 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 115.2550 0.0000 115.3450 0.4700 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 112.2550 0.0000 112.3450 0.4700 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 109.2550 0.0000 109.3450 0.4700 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 106.2550 0.0000 106.3450 0.4700 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 103.2550 0.0000 103.3450 0.4700 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 100.2550 0.0000 100.3450 0.4700 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 97.2550 0.0000 97.3450 0.4700 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 94.2550 0.0000 94.3450 0.4700 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 91.2550 0.0000 91.3450 0.4700 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 88.2550 0.0000 88.3450 0.4700 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 85.2550 0.0000 85.3450 0.4700 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 82.2550 0.0000 82.3450 0.4700 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 79.2550 0.0000 79.3450 0.4700 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 76.2550 0.0000 76.3450 0.4700 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 73.2550 0.0000 73.3450 0.4700 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 70.2550 0.0000 70.3450 0.4700 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 67.2550 0.0000 67.3450 0.4700 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 64.2550 0.0000 64.3450 0.4700 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 61.2550 0.0000 61.3450 0.4700 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 58.2550 0.0000 58.3450 0.4700 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 55.2550 0.0000 55.3450 0.4700 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 52.2550 0.0000 52.3450 0.4700 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 49.2550 0.0000 49.3450 0.4700 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 46.2550 0.0000 46.3450 0.4700 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 43.2550 0.0000 43.3450 0.4700 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 40.2550 0.0000 40.3450 0.4700 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 37.2550 0.0000 37.3450 0.4700 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 34.2550 0.0000 34.3450 0.4700 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 31.2550 0.0000 31.3450 0.4700 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 28.2550 0.0000 28.3450 0.4700 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 25.2550 0.0000 25.3450 0.4700 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 22.2550 0.0000 22.3450 0.4700 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 19.2550 0.0000 19.3450 0.4700 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 16.2550 0.0000 16.3450 0.4700 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.2550 0.0000 13.3450 0.4700 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.2550 0.0000 10.3450 0.4700 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 164.7500 0.5200 164.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 159.7500 0.5200 159.8500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 154.7500 0.5200 154.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 149.7500 0.5200 149.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 144.7500 0.5200 144.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 139.7500 0.5200 139.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 134.7500 0.5200 134.8500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 129.7500 0.5200 129.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 124.7500 0.5200 124.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 119.7500 0.5200 119.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 114.7500 0.5200 114.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 109.7500 0.5200 109.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 104.7500 0.5200 104.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 99.7500 0.5200 99.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 94.7500 0.5200 94.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 89.7500 0.5200 89.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 84.7500 0.5200 84.8500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 287.2550 569.5300 287.3450 570.0000 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 287.5050 569.3700 570.0000 570.0000 ;
      RECT 282.5050 569.3700 287.0950 570.0000 ;
      RECT 0.0000 569.3700 282.0950 570.0000 ;
      RECT 0.0000 0.6300 570.0000 569.3700 ;
      RECT 559.5050 0.0000 570.0000 0.6300 ;
      RECT 556.5050 0.0000 559.0950 0.6300 ;
      RECT 553.5050 0.0000 556.0950 0.6300 ;
      RECT 550.5050 0.0000 553.0950 0.6300 ;
      RECT 547.5050 0.0000 550.0950 0.6300 ;
      RECT 544.5050 0.0000 547.0950 0.6300 ;
      RECT 541.5050 0.0000 544.0950 0.6300 ;
      RECT 538.5050 0.0000 541.0950 0.6300 ;
      RECT 535.5050 0.0000 538.0950 0.6300 ;
      RECT 532.5050 0.0000 535.0950 0.6300 ;
      RECT 529.5050 0.0000 532.0950 0.6300 ;
      RECT 526.5050 0.0000 529.0950 0.6300 ;
      RECT 523.5050 0.0000 526.0950 0.6300 ;
      RECT 520.5050 0.0000 523.0950 0.6300 ;
      RECT 517.5050 0.0000 520.0950 0.6300 ;
      RECT 514.5050 0.0000 517.0950 0.6300 ;
      RECT 511.5050 0.0000 514.0950 0.6300 ;
      RECT 508.5050 0.0000 511.0950 0.6300 ;
      RECT 505.5050 0.0000 508.0950 0.6300 ;
      RECT 502.5050 0.0000 505.0950 0.6300 ;
      RECT 499.5050 0.0000 502.0950 0.6300 ;
      RECT 496.5050 0.0000 499.0950 0.6300 ;
      RECT 493.5050 0.0000 496.0950 0.6300 ;
      RECT 490.5050 0.0000 493.0950 0.6300 ;
      RECT 487.5050 0.0000 490.0950 0.6300 ;
      RECT 484.5050 0.0000 487.0950 0.6300 ;
      RECT 481.5050 0.0000 484.0950 0.6300 ;
      RECT 478.5050 0.0000 481.0950 0.6300 ;
      RECT 475.5050 0.0000 478.0950 0.6300 ;
      RECT 472.5050 0.0000 475.0950 0.6300 ;
      RECT 469.5050 0.0000 472.0950 0.6300 ;
      RECT 466.5050 0.0000 469.0950 0.6300 ;
      RECT 463.5050 0.0000 466.0950 0.6300 ;
      RECT 460.5050 0.0000 463.0950 0.6300 ;
      RECT 457.5050 0.0000 460.0950 0.6300 ;
      RECT 454.5050 0.0000 457.0950 0.6300 ;
      RECT 451.5050 0.0000 454.0950 0.6300 ;
      RECT 448.5050 0.0000 451.0950 0.6300 ;
      RECT 445.5050 0.0000 448.0950 0.6300 ;
      RECT 442.5050 0.0000 445.0950 0.6300 ;
      RECT 439.5050 0.0000 442.0950 0.6300 ;
      RECT 436.5050 0.0000 439.0950 0.6300 ;
      RECT 433.5050 0.0000 436.0950 0.6300 ;
      RECT 430.5050 0.0000 433.0950 0.6300 ;
      RECT 427.5050 0.0000 430.0950 0.6300 ;
      RECT 424.5050 0.0000 427.0950 0.6300 ;
      RECT 421.5050 0.0000 424.0950 0.6300 ;
      RECT 418.5050 0.0000 421.0950 0.6300 ;
      RECT 415.5050 0.0000 418.0950 0.6300 ;
      RECT 412.5050 0.0000 415.0950 0.6300 ;
      RECT 409.5050 0.0000 412.0950 0.6300 ;
      RECT 406.5050 0.0000 409.0950 0.6300 ;
      RECT 403.5050 0.0000 406.0950 0.6300 ;
      RECT 400.5050 0.0000 403.0950 0.6300 ;
      RECT 397.5050 0.0000 400.0950 0.6300 ;
      RECT 394.5050 0.0000 397.0950 0.6300 ;
      RECT 391.5050 0.0000 394.0950 0.6300 ;
      RECT 388.5050 0.0000 391.0950 0.6300 ;
      RECT 385.5050 0.0000 388.0950 0.6300 ;
      RECT 382.5050 0.0000 385.0950 0.6300 ;
      RECT 379.5050 0.0000 382.0950 0.6300 ;
      RECT 376.5050 0.0000 379.0950 0.6300 ;
      RECT 373.5050 0.0000 376.0950 0.6300 ;
      RECT 370.5050 0.0000 373.0950 0.6300 ;
      RECT 367.5050 0.0000 370.0950 0.6300 ;
      RECT 364.5050 0.0000 367.0950 0.6300 ;
      RECT 361.5050 0.0000 364.0950 0.6300 ;
      RECT 358.5050 0.0000 361.0950 0.6300 ;
      RECT 355.5050 0.0000 358.0950 0.6300 ;
      RECT 352.5050 0.0000 355.0950 0.6300 ;
      RECT 349.5050 0.0000 352.0950 0.6300 ;
      RECT 346.5050 0.0000 349.0950 0.6300 ;
      RECT 343.5050 0.0000 346.0950 0.6300 ;
      RECT 340.5050 0.0000 343.0950 0.6300 ;
      RECT 337.5050 0.0000 340.0950 0.6300 ;
      RECT 334.5050 0.0000 337.0950 0.6300 ;
      RECT 331.5050 0.0000 334.0950 0.6300 ;
      RECT 328.5050 0.0000 331.0950 0.6300 ;
      RECT 325.5050 0.0000 328.0950 0.6300 ;
      RECT 322.5050 0.0000 325.0950 0.6300 ;
      RECT 319.5050 0.0000 322.0950 0.6300 ;
      RECT 316.5050 0.0000 319.0950 0.6300 ;
      RECT 313.5050 0.0000 316.0950 0.6300 ;
      RECT 310.5050 0.0000 313.0950 0.6300 ;
      RECT 307.5050 0.0000 310.0950 0.6300 ;
      RECT 304.5050 0.0000 307.0950 0.6300 ;
      RECT 301.5050 0.0000 304.0950 0.6300 ;
      RECT 298.5050 0.0000 301.0950 0.6300 ;
      RECT 295.5050 0.0000 298.0950 0.6300 ;
      RECT 292.5050 0.0000 295.0950 0.6300 ;
      RECT 289.5050 0.0000 292.0950 0.6300 ;
      RECT 286.5050 0.0000 289.0950 0.6300 ;
      RECT 283.5050 0.0000 286.0950 0.6300 ;
      RECT 280.5050 0.0000 283.0950 0.6300 ;
      RECT 277.5050 0.0000 280.0950 0.6300 ;
      RECT 274.5050 0.0000 277.0950 0.6300 ;
      RECT 271.5050 0.0000 274.0950 0.6300 ;
      RECT 268.5050 0.0000 271.0950 0.6300 ;
      RECT 265.5050 0.0000 268.0950 0.6300 ;
      RECT 262.5050 0.0000 265.0950 0.6300 ;
      RECT 259.5050 0.0000 262.0950 0.6300 ;
      RECT 256.5050 0.0000 259.0950 0.6300 ;
      RECT 253.5050 0.0000 256.0950 0.6300 ;
      RECT 250.5050 0.0000 253.0950 0.6300 ;
      RECT 247.5050 0.0000 250.0950 0.6300 ;
      RECT 244.5050 0.0000 247.0950 0.6300 ;
      RECT 241.5050 0.0000 244.0950 0.6300 ;
      RECT 238.5050 0.0000 241.0950 0.6300 ;
      RECT 235.5050 0.0000 238.0950 0.6300 ;
      RECT 232.5050 0.0000 235.0950 0.6300 ;
      RECT 229.5050 0.0000 232.0950 0.6300 ;
      RECT 226.5050 0.0000 229.0950 0.6300 ;
      RECT 223.5050 0.0000 226.0950 0.6300 ;
      RECT 220.5050 0.0000 223.0950 0.6300 ;
      RECT 217.5050 0.0000 220.0950 0.6300 ;
      RECT 214.5050 0.0000 217.0950 0.6300 ;
      RECT 211.5050 0.0000 214.0950 0.6300 ;
      RECT 208.5050 0.0000 211.0950 0.6300 ;
      RECT 205.5050 0.0000 208.0950 0.6300 ;
      RECT 202.5050 0.0000 205.0950 0.6300 ;
      RECT 199.5050 0.0000 202.0950 0.6300 ;
      RECT 196.5050 0.0000 199.0950 0.6300 ;
      RECT 193.5050 0.0000 196.0950 0.6300 ;
      RECT 190.5050 0.0000 193.0950 0.6300 ;
      RECT 187.5050 0.0000 190.0950 0.6300 ;
      RECT 184.5050 0.0000 187.0950 0.6300 ;
      RECT 181.5050 0.0000 184.0950 0.6300 ;
      RECT 178.5050 0.0000 181.0950 0.6300 ;
      RECT 175.5050 0.0000 178.0950 0.6300 ;
      RECT 172.5050 0.0000 175.0950 0.6300 ;
      RECT 169.5050 0.0000 172.0950 0.6300 ;
      RECT 166.5050 0.0000 169.0950 0.6300 ;
      RECT 163.5050 0.0000 166.0950 0.6300 ;
      RECT 160.5050 0.0000 163.0950 0.6300 ;
      RECT 157.5050 0.0000 160.0950 0.6300 ;
      RECT 154.5050 0.0000 157.0950 0.6300 ;
      RECT 151.5050 0.0000 154.0950 0.6300 ;
      RECT 148.5050 0.0000 151.0950 0.6300 ;
      RECT 145.5050 0.0000 148.0950 0.6300 ;
      RECT 142.5050 0.0000 145.0950 0.6300 ;
      RECT 139.5050 0.0000 142.0950 0.6300 ;
      RECT 136.5050 0.0000 139.0950 0.6300 ;
      RECT 133.5050 0.0000 136.0950 0.6300 ;
      RECT 130.5050 0.0000 133.0950 0.6300 ;
      RECT 127.5050 0.0000 130.0950 0.6300 ;
      RECT 124.5050 0.0000 127.0950 0.6300 ;
      RECT 121.5050 0.0000 124.0950 0.6300 ;
      RECT 118.5050 0.0000 121.0950 0.6300 ;
      RECT 115.5050 0.0000 118.0950 0.6300 ;
      RECT 112.5050 0.0000 115.0950 0.6300 ;
      RECT 109.5050 0.0000 112.0950 0.6300 ;
      RECT 106.5050 0.0000 109.0950 0.6300 ;
      RECT 103.5050 0.0000 106.0950 0.6300 ;
      RECT 100.5050 0.0000 103.0950 0.6300 ;
      RECT 97.5050 0.0000 100.0950 0.6300 ;
      RECT 94.5050 0.0000 97.0950 0.6300 ;
      RECT 91.5050 0.0000 94.0950 0.6300 ;
      RECT 88.5050 0.0000 91.0950 0.6300 ;
      RECT 85.5050 0.0000 88.0950 0.6300 ;
      RECT 82.5050 0.0000 85.0950 0.6300 ;
      RECT 79.5050 0.0000 82.0950 0.6300 ;
      RECT 76.5050 0.0000 79.0950 0.6300 ;
      RECT 73.5050 0.0000 76.0950 0.6300 ;
      RECT 70.5050 0.0000 73.0950 0.6300 ;
      RECT 67.5050 0.0000 70.0950 0.6300 ;
      RECT 64.5050 0.0000 67.0950 0.6300 ;
      RECT 61.5050 0.0000 64.0950 0.6300 ;
      RECT 58.5050 0.0000 61.0950 0.6300 ;
      RECT 55.5050 0.0000 58.0950 0.6300 ;
      RECT 52.5050 0.0000 55.0950 0.6300 ;
      RECT 49.5050 0.0000 52.0950 0.6300 ;
      RECT 46.5050 0.0000 49.0950 0.6300 ;
      RECT 43.5050 0.0000 46.0950 0.6300 ;
      RECT 40.5050 0.0000 43.0950 0.6300 ;
      RECT 37.5050 0.0000 40.0950 0.6300 ;
      RECT 34.5050 0.0000 37.0950 0.6300 ;
      RECT 31.5050 0.0000 34.0950 0.6300 ;
      RECT 28.5050 0.0000 31.0950 0.6300 ;
      RECT 25.5050 0.0000 28.0950 0.6300 ;
      RECT 22.5050 0.0000 25.0950 0.6300 ;
      RECT 19.5050 0.0000 22.0950 0.6300 ;
      RECT 16.5050 0.0000 19.0950 0.6300 ;
      RECT 13.5050 0.0000 16.0950 0.6300 ;
      RECT 10.5050 0.0000 13.0950 0.6300 ;
      RECT 0.0000 0.0000 10.0950 0.6300 ;
    LAYER M2 ;
      RECT 0.0000 485.0100 570.0000 570.0000 ;
      RECT 0.6800 484.5900 570.0000 485.0100 ;
      RECT 0.0000 480.0100 570.0000 484.5900 ;
      RECT 0.6800 479.5900 570.0000 480.0100 ;
      RECT 0.0000 475.0100 570.0000 479.5900 ;
      RECT 0.6800 474.5900 570.0000 475.0100 ;
      RECT 0.0000 470.0100 570.0000 474.5900 ;
      RECT 0.6800 469.5900 570.0000 470.0100 ;
      RECT 0.0000 465.0100 570.0000 469.5900 ;
      RECT 0.6800 464.5900 570.0000 465.0100 ;
      RECT 0.0000 460.0100 570.0000 464.5900 ;
      RECT 0.6800 459.5900 570.0000 460.0100 ;
      RECT 0.0000 455.0100 570.0000 459.5900 ;
      RECT 0.6800 454.5900 570.0000 455.0100 ;
      RECT 0.0000 450.0100 570.0000 454.5900 ;
      RECT 0.6800 449.5900 570.0000 450.0100 ;
      RECT 0.0000 445.0100 570.0000 449.5900 ;
      RECT 0.6800 444.5900 570.0000 445.0100 ;
      RECT 0.0000 440.0100 570.0000 444.5900 ;
      RECT 0.6800 439.5900 570.0000 440.0100 ;
      RECT 0.0000 435.0100 570.0000 439.5900 ;
      RECT 0.6800 434.5900 570.0000 435.0100 ;
      RECT 0.0000 430.0100 570.0000 434.5900 ;
      RECT 0.6800 429.5900 570.0000 430.0100 ;
      RECT 0.0000 425.0100 570.0000 429.5900 ;
      RECT 0.6800 424.5900 570.0000 425.0100 ;
      RECT 0.0000 420.0100 570.0000 424.5900 ;
      RECT 0.6800 419.5900 570.0000 420.0100 ;
      RECT 0.0000 415.0100 570.0000 419.5900 ;
      RECT 0.6800 414.5900 570.0000 415.0100 ;
      RECT 0.0000 410.0100 570.0000 414.5900 ;
      RECT 0.6800 409.5900 570.0000 410.0100 ;
      RECT 0.0000 405.0100 570.0000 409.5900 ;
      RECT 0.6800 404.5900 570.0000 405.0100 ;
      RECT 0.0000 400.0100 570.0000 404.5900 ;
      RECT 0.6800 399.5900 570.0000 400.0100 ;
      RECT 0.0000 395.0100 570.0000 399.5900 ;
      RECT 0.6800 394.5900 570.0000 395.0100 ;
      RECT 0.0000 390.0100 570.0000 394.5900 ;
      RECT 0.6800 389.5900 570.0000 390.0100 ;
      RECT 0.0000 385.0100 570.0000 389.5900 ;
      RECT 0.6800 384.5900 570.0000 385.0100 ;
      RECT 0.0000 380.0100 570.0000 384.5900 ;
      RECT 0.6800 379.5900 570.0000 380.0100 ;
      RECT 0.0000 375.0100 570.0000 379.5900 ;
      RECT 0.6800 374.5900 570.0000 375.0100 ;
      RECT 0.0000 370.0100 570.0000 374.5900 ;
      RECT 0.6800 369.5900 570.0000 370.0100 ;
      RECT 0.0000 365.0100 570.0000 369.5900 ;
      RECT 0.6800 364.5900 570.0000 365.0100 ;
      RECT 0.0000 360.0100 570.0000 364.5900 ;
      RECT 0.6800 359.5900 570.0000 360.0100 ;
      RECT 0.0000 355.0100 570.0000 359.5900 ;
      RECT 0.6800 354.5900 570.0000 355.0100 ;
      RECT 0.0000 350.0100 570.0000 354.5900 ;
      RECT 0.6800 349.5900 570.0000 350.0100 ;
      RECT 0.0000 345.0100 570.0000 349.5900 ;
      RECT 0.6800 344.5900 570.0000 345.0100 ;
      RECT 0.0000 340.0100 570.0000 344.5900 ;
      RECT 0.6800 339.5900 570.0000 340.0100 ;
      RECT 0.0000 335.0100 570.0000 339.5900 ;
      RECT 0.6800 334.5900 570.0000 335.0100 ;
      RECT 0.0000 330.0100 570.0000 334.5900 ;
      RECT 0.6800 329.5900 570.0000 330.0100 ;
      RECT 0.0000 325.0100 570.0000 329.5900 ;
      RECT 0.6800 324.5900 570.0000 325.0100 ;
      RECT 0.0000 320.0100 570.0000 324.5900 ;
      RECT 0.6800 319.5900 570.0000 320.0100 ;
      RECT 0.0000 315.0100 570.0000 319.5900 ;
      RECT 0.6800 314.5900 570.0000 315.0100 ;
      RECT 0.0000 310.0100 570.0000 314.5900 ;
      RECT 0.6800 309.5900 570.0000 310.0100 ;
      RECT 0.0000 305.0100 570.0000 309.5900 ;
      RECT 0.6800 304.5900 570.0000 305.0100 ;
      RECT 0.0000 300.0100 570.0000 304.5900 ;
      RECT 0.6800 299.5900 570.0000 300.0100 ;
      RECT 0.0000 295.0100 570.0000 299.5900 ;
      RECT 0.6800 294.5900 570.0000 295.0100 ;
      RECT 0.0000 290.0100 570.0000 294.5900 ;
      RECT 0.6800 289.5900 570.0000 290.0100 ;
      RECT 0.0000 285.0100 570.0000 289.5900 ;
      RECT 0.6800 284.5900 570.0000 285.0100 ;
      RECT 0.0000 280.0100 570.0000 284.5900 ;
      RECT 0.6800 279.5900 570.0000 280.0100 ;
      RECT 0.0000 275.0100 570.0000 279.5900 ;
      RECT 0.6800 274.5900 570.0000 275.0100 ;
      RECT 0.0000 270.0100 570.0000 274.5900 ;
      RECT 0.6800 269.5900 570.0000 270.0100 ;
      RECT 0.0000 265.0100 570.0000 269.5900 ;
      RECT 0.6800 264.5900 570.0000 265.0100 ;
      RECT 0.0000 260.0100 570.0000 264.5900 ;
      RECT 0.6800 259.5900 570.0000 260.0100 ;
      RECT 0.0000 255.0100 570.0000 259.5900 ;
      RECT 0.6800 254.5900 570.0000 255.0100 ;
      RECT 0.0000 250.0100 570.0000 254.5900 ;
      RECT 0.6800 249.5900 570.0000 250.0100 ;
      RECT 0.0000 245.0100 570.0000 249.5900 ;
      RECT 0.6800 244.5900 570.0000 245.0100 ;
      RECT 0.0000 240.0100 570.0000 244.5900 ;
      RECT 0.6800 239.5900 570.0000 240.0100 ;
      RECT 0.0000 235.0100 570.0000 239.5900 ;
      RECT 0.6800 234.5900 570.0000 235.0100 ;
      RECT 0.0000 230.0100 570.0000 234.5900 ;
      RECT 0.6800 229.5900 570.0000 230.0100 ;
      RECT 0.0000 225.0100 570.0000 229.5900 ;
      RECT 0.6800 224.5900 570.0000 225.0100 ;
      RECT 0.0000 220.0100 570.0000 224.5900 ;
      RECT 0.6800 219.5900 570.0000 220.0100 ;
      RECT 0.0000 215.0100 570.0000 219.5900 ;
      RECT 0.6800 214.5900 570.0000 215.0100 ;
      RECT 0.0000 210.0100 570.0000 214.5900 ;
      RECT 0.6800 209.5900 570.0000 210.0100 ;
      RECT 0.0000 205.0100 570.0000 209.5900 ;
      RECT 0.6800 204.5900 570.0000 205.0100 ;
      RECT 0.0000 200.0100 570.0000 204.5900 ;
      RECT 0.6800 199.5900 570.0000 200.0100 ;
      RECT 0.0000 195.0100 570.0000 199.5900 ;
      RECT 0.6800 194.5900 570.0000 195.0100 ;
      RECT 0.0000 190.0100 570.0000 194.5900 ;
      RECT 0.6800 189.5900 570.0000 190.0100 ;
      RECT 0.0000 185.0100 570.0000 189.5900 ;
      RECT 0.6800 184.5900 570.0000 185.0100 ;
      RECT 0.0000 180.0100 570.0000 184.5900 ;
      RECT 0.6800 179.5900 570.0000 180.0100 ;
      RECT 0.0000 175.0100 570.0000 179.5900 ;
      RECT 0.6800 174.5900 570.0000 175.0100 ;
      RECT 0.0000 170.0100 570.0000 174.5900 ;
      RECT 0.6800 169.5900 570.0000 170.0100 ;
      RECT 0.0000 165.0100 570.0000 169.5900 ;
      RECT 0.6800 164.5900 570.0000 165.0100 ;
      RECT 0.0000 160.0100 570.0000 164.5900 ;
      RECT 0.6800 159.5900 570.0000 160.0100 ;
      RECT 0.0000 155.0100 570.0000 159.5900 ;
      RECT 0.6800 154.5900 570.0000 155.0100 ;
      RECT 0.0000 150.0100 570.0000 154.5900 ;
      RECT 0.6800 149.5900 570.0000 150.0100 ;
      RECT 0.0000 145.0100 570.0000 149.5900 ;
      RECT 0.6800 144.5900 570.0000 145.0100 ;
      RECT 0.0000 140.0100 570.0000 144.5900 ;
      RECT 0.6800 139.5900 570.0000 140.0100 ;
      RECT 0.0000 135.0100 570.0000 139.5900 ;
      RECT 0.6800 134.5900 570.0000 135.0100 ;
      RECT 0.0000 130.0100 570.0000 134.5900 ;
      RECT 0.6800 129.5900 570.0000 130.0100 ;
      RECT 0.0000 125.0100 570.0000 129.5900 ;
      RECT 0.6800 124.5900 570.0000 125.0100 ;
      RECT 0.0000 120.0100 570.0000 124.5900 ;
      RECT 0.6800 119.5900 570.0000 120.0100 ;
      RECT 0.0000 115.0100 570.0000 119.5900 ;
      RECT 0.6800 114.5900 570.0000 115.0100 ;
      RECT 0.0000 110.0100 570.0000 114.5900 ;
      RECT 0.6800 109.5900 570.0000 110.0100 ;
      RECT 0.0000 105.0100 570.0000 109.5900 ;
      RECT 0.6800 104.5900 570.0000 105.0100 ;
      RECT 0.0000 100.0100 570.0000 104.5900 ;
      RECT 0.6800 99.5900 570.0000 100.0100 ;
      RECT 0.0000 95.0100 570.0000 99.5900 ;
      RECT 0.6800 94.5900 570.0000 95.0100 ;
      RECT 0.0000 90.0100 570.0000 94.5900 ;
      RECT 0.6800 89.5900 570.0000 90.0100 ;
      RECT 0.0000 85.0100 570.0000 89.5900 ;
      RECT 0.6800 84.5900 570.0000 85.0100 ;
      RECT 0.0000 0.0000 570.0000 84.5900 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 570.0000 570.0000 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 570.0000 570.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 570.0000 570.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 570.0000 570.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 570.0000 570.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 570.0000 570.0000 ;
  END
END core

END LIBRARY
